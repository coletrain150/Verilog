library verilog;
use verilog.vl_types.all;
entity tb_sync is
end tb_sync;
