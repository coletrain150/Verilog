library verilog;
use verilog.vl_types.all;
entity flex_counter_NUM_CNT_BITS8_ROLLOVER_VAL9_DW01_inc_1 is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        SUM             : out    vl_logic_vector(7 downto 0)
    );
end flex_counter_NUM_CNT_BITS8_ROLLOVER_VAL9_DW01_inc_1;
