// $Id: $
// File name:   tb_decode.sv
// Created:     3/10/2014
// Author:      Cole Reinhold
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: decoder test bench
// ,
