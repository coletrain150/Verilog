
module sync ( clk, n_reset, async_in, sync_out );
  input clk, n_reset, async_in;
  output sync_out;
  wire   out_one;

  DFFSR out_one_reg ( .D(async_in), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        out_one) );
  DFFSR sec_out_reg ( .D(out_one), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        sync_out) );
endmodule


module controller ( clk, n_reset, dr, overflow, cnt_up, modwait, op, src1, 
        src2, dest, err );
  output [1:0] op;
  output [3:0] src1;
  output [3:0] src2;
  output [3:0] dest;
  input clk, n_reset, dr, overflow;
  output cnt_up, modwait, err;
  wire   nextflag, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76;
  wire   [3:0] state;
  wire   [3:0] nextstate;
  assign dest[3] = 1'b0;
  assign src2[3] = 1'b0;
  assign src1[3] = 1'b0;

  DFFSR \state_reg[0]  ( .D(nextstate[0]), .CLK(clk), .R(n_reset), .S(1'b1), 
        .Q(state[0]) );
  DFFSR \state_reg[2]  ( .D(nextstate[2]), .CLK(clk), .R(n_reset), .S(1'b1), 
        .Q(state[2]) );
  DFFSR \state_reg[1]  ( .D(nextstate[1]), .CLK(clk), .R(n_reset), .S(1'b1), 
        .Q(state[1]) );
  DFFSR \state_reg[3]  ( .D(nextstate[3]), .CLK(clk), .R(n_reset), .S(1'b1), 
        .Q(state[3]) );
  DFFSR flag_reg ( .D(nextflag), .CLK(clk), .R(n_reset), .S(1'b1), .Q(modwait)
         );
  INVX4 U8 ( .A(n29), .Y(n22) );
  BUFX2 U9 ( .A(state[2]), .Y(n6) );
  INVX2 U10 ( .A(n22), .Y(n23) );
  INVX2 U11 ( .A(n9), .Y(n16) );
  INVX2 U12 ( .A(n9), .Y(n18) );
  INVX2 U13 ( .A(overflow), .Y(n7) );
  INVX2 U14 ( .A(overflow), .Y(n55) );
  BUFX2 U15 ( .A(n55), .Y(n8) );
  INVX1 U16 ( .A(n53), .Y(n43) );
  INVX1 U17 ( .A(n48), .Y(n49) );
  INVX1 U18 ( .A(n48), .Y(n45) );
  BUFX4 U19 ( .A(state[1]), .Y(n9) );
  BUFX2 U20 ( .A(state[1]), .Y(n21) );
  INVX2 U21 ( .A(n14), .Y(n10) );
  BUFX2 U22 ( .A(n62), .Y(n11) );
  INVX1 U23 ( .A(op[0]), .Y(n73) );
  BUFX4 U24 ( .A(n34), .Y(n12) );
  BUFX2 U25 ( .A(n74), .Y(n13) );
  INVX1 U26 ( .A(state[0]), .Y(n74) );
  INVX1 U27 ( .A(src1[2]), .Y(n14) );
  INVX2 U28 ( .A(n60), .Y(src1[2]) );
  BUFX2 U29 ( .A(n68), .Y(n15) );
  INVX1 U30 ( .A(n63), .Y(n17) );
  INVX1 U31 ( .A(src2[0]), .Y(n19) );
  INVX2 U32 ( .A(n19), .Y(n20) );
  INVX4 U33 ( .A(n37), .Y(n63) );
  BUFX2 U34 ( .A(src2[1]), .Y(n24) );
  INVX2 U35 ( .A(n26), .Y(n25) );
  INVX1 U36 ( .A(src1[1]), .Y(n26) );
  INVX1 U37 ( .A(n30), .Y(n27) );
  INVX2 U38 ( .A(n18), .Y(n30) );
  BUFX2 U39 ( .A(n61), .Y(n28) );
  BUFX2 U40 ( .A(state[2]), .Y(n29) );
  OR2X2 U41 ( .A(n6), .B(n21), .Y(n61) );
  AND2X2 U42 ( .A(n29), .B(n21), .Y(n31) );
  INVX1 U43 ( .A(n31), .Y(n51) );
  AND2X2 U44 ( .A(n34), .B(n35), .Y(n32) );
  INVX1 U45 ( .A(n32), .Y(n69) );
  INVX2 U46 ( .A(n37), .Y(n70) );
  NAND3X1 U47 ( .A(n6), .B(n9), .C(n63), .Y(n33) );
  OR2X2 U48 ( .A(n28), .B(n11), .Y(n68) );
  AND2X2 U49 ( .A(n22), .B(n18), .Y(n34) );
  INVX4 U50 ( .A(n66), .Y(src1[0]) );
  BUFX4 U51 ( .A(state[0]), .Y(n35) );
  AND2X1 U52 ( .A(n68), .B(n67), .Y(n72) );
  INVX4 U53 ( .A(n38), .Y(src2[2]) );
  INVX4 U54 ( .A(n52), .Y(src2[0]) );
  INVX4 U55 ( .A(n33), .Y(src2[1]) );
  INVX2 U56 ( .A(state[3]), .Y(n36) );
  INVX4 U57 ( .A(n36), .Y(n37) );
  OR2X2 U58 ( .A(n61), .B(n62), .Y(n38) );
  INVX4 U59 ( .A(n59), .Y(src1[1]) );
  NAND3X1 U60 ( .A(n30), .B(n70), .C(n23), .Y(n67) );
  OAI22X1 U61 ( .A(n67), .B(n7), .C(dr), .D(n69), .Y(n53) );
  NAND2X1 U62 ( .A(n32), .B(n17), .Y(n56) );
  NOR2X1 U63 ( .A(n70), .B(n55), .Y(n41) );
  NAND2X1 U64 ( .A(n51), .B(n70), .Y(n75) );
  INVX2 U65 ( .A(n75), .Y(n58) );
  AOI21X1 U66 ( .A(dr), .B(n58), .C(n24), .Y(n39) );
  OAI21X1 U67 ( .A(n12), .B(n75), .C(n39), .Y(n40) );
  AOI22X1 U68 ( .A(n41), .B(n12), .C(n40), .D(n13), .Y(n42) );
  NAND3X1 U69 ( .A(n56), .B(n43), .C(n42), .Y(nextstate[0]) );
  NAND3X1 U70 ( .A(n35), .B(n27), .C(n70), .Y(n44) );
  INVX2 U71 ( .A(n44), .Y(dest[2]) );
  OAI21X1 U72 ( .A(dr), .B(n23), .C(dest[2]), .Y(n47) );
  NAND3X1 U73 ( .A(n70), .B(n13), .C(n55), .Y(n48) );
  NAND2X1 U74 ( .A(n45), .B(n30), .Y(n46) );
  NAND3X1 U75 ( .A(n63), .B(n9), .C(n22), .Y(n59) );
  NAND2X1 U76 ( .A(n25), .B(n13), .Y(n76) );
  NAND3X1 U77 ( .A(n47), .B(n76), .C(n46), .Y(nextstate[1]) );
  NAND3X1 U78 ( .A(n6), .B(n63), .C(n16), .Y(n60) );
  AOI21X1 U79 ( .A(n49), .B(n23), .C(n10), .Y(n50) );
  OAI21X1 U80 ( .A(n26), .B(n13), .C(n50), .Y(nextstate[2]) );
  NAND2X1 U81 ( .A(n37), .B(n74), .Y(n62) );
  NAND3X1 U82 ( .A(n35), .B(n70), .C(n31), .Y(n52) );
  NOR2X1 U83 ( .A(n20), .B(n53), .Y(n54) );
  OAI21X1 U84 ( .A(n8), .B(n15), .C(n54), .Y(nextstate[3]) );
  INVX2 U85 ( .A(n56), .Y(err) );
  OAI21X1 U86 ( .A(n35), .B(n12), .C(n69), .Y(n57) );
  AND2X2 U87 ( .A(n58), .B(n57), .Y(dest[0]) );
  MUX2X1 U88 ( .B(n14), .A(n26), .S(n35), .Y(dest[1]) );
  OAI21X1 U89 ( .A(n16), .B(n22), .C(n63), .Y(n64) );
  AOI22X1 U90 ( .A(n35), .B(n64), .C(n22), .D(n18), .Y(n65) );
  OAI21X1 U91 ( .A(src2[1]), .B(n35), .C(n65), .Y(n66) );
  OAI21X1 U92 ( .A(n17), .B(n12), .C(n68), .Y(op[0]) );
  NAND2X1 U93 ( .A(n32), .B(n70), .Y(n71) );
  NAND2X1 U94 ( .A(n71), .B(n72), .Y(op[1]) );
  OAI21X1 U95 ( .A(n75), .B(n13), .C(n73), .Y(nextflag) );
  INVX2 U96 ( .A(n76), .Y(cnt_up) );
endmodule


module datapath_ctrl ( op, w_data_sel, w_en, alu_op );
  input [1:0] op;
  output w_data_sel, w_en, alu_op;
  wire   \op[0] , n1, n2;
  assign w_data_sel = \op[0] ;
  assign \op[0]  = op[0];

  AND2X2 U1 ( .A(op[1]), .B(\op[0] ), .Y(alu_op) );
  INVX1 U2 ( .A(op[1]), .Y(n1) );
  INVX1 U3 ( .A(\op[0] ), .Y(n2) );
  NAND2X1 U4 ( .A(n2), .B(n1), .Y(w_en) );
endmodule


module regfile_NUM_REG_ADDR_BITS4_REG_SIZE_BITS16 ( clk, n_reset, w_sel, 
        r1_sel, r2_sel, w_data, w_en, r1_data, r2_data, outreg_data );
  input [3:0] w_sel;
  input [3:0] r1_sel;
  input [3:0] r2_sel;
  input [15:0] w_data;
  output [15:0] r1_data;
  output [15:0] r2_data;
  output [15:0] outreg_data;
  input clk, n_reset, w_en;
  wire   \regs[15][15] , \regs[15][14] , \regs[15][13] , \regs[15][12] ,
         \regs[15][11] , \regs[15][10] , \regs[15][9] , \regs[15][8] ,
         \regs[15][7] , \regs[15][6] , \regs[15][5] , \regs[15][4] ,
         \regs[15][3] , \regs[15][2] , \regs[15][1] , \regs[15][0] ,
         \regs[14][15] , \regs[14][14] , \regs[14][13] , \regs[14][12] ,
         \regs[14][11] , \regs[14][10] , \regs[14][9] , \regs[14][8] ,
         \regs[14][7] , \regs[14][6] , \regs[14][5] , \regs[14][4] ,
         \regs[14][3] , \regs[14][2] , \regs[14][1] , \regs[14][0] ,
         \regs[13][15] , \regs[13][14] , \regs[13][13] , \regs[13][12] ,
         \regs[13][11] , \regs[13][10] , \regs[13][9] , \regs[13][8] ,
         \regs[13][7] , \regs[13][6] , \regs[13][5] , \regs[13][4] ,
         \regs[13][3] , \regs[13][2] , \regs[13][1] , \regs[13][0] ,
         \regs[12][15] , \regs[12][14] , \regs[12][13] , \regs[12][12] ,
         \regs[12][11] , \regs[12][10] , \regs[12][9] , \regs[12][8] ,
         \regs[12][7] , \regs[12][6] , \regs[12][5] , \regs[12][4] ,
         \regs[12][3] , \regs[12][2] , \regs[12][1] , \regs[12][0] ,
         \regs[11][15] , \regs[11][14] , \regs[11][13] , \regs[11][12] ,
         \regs[11][11] , \regs[11][10] , \regs[11][9] , \regs[11][8] ,
         \regs[11][7] , \regs[11][6] , \regs[11][5] , \regs[11][4] ,
         \regs[11][3] , \regs[11][2] , \regs[11][1] , \regs[11][0] ,
         \regs[10][15] , \regs[10][14] , \regs[10][13] , \regs[10][12] ,
         \regs[10][11] , \regs[10][10] , \regs[10][9] , \regs[10][8] ,
         \regs[10][7] , \regs[10][6] , \regs[10][5] , \regs[10][4] ,
         \regs[10][3] , \regs[10][2] , \regs[10][1] , \regs[10][0] ,
         \regs[9][15] , \regs[9][14] , \regs[9][13] , \regs[9][12] ,
         \regs[9][11] , \regs[9][10] , \regs[9][9] , \regs[9][8] ,
         \regs[9][7] , \regs[9][6] , \regs[9][5] , \regs[9][4] , \regs[9][3] ,
         \regs[9][2] , \regs[9][1] , \regs[9][0] , \regs[8][15] ,
         \regs[8][14] , \regs[8][13] , \regs[8][12] , \regs[8][11] ,
         \regs[8][10] , \regs[8][9] , \regs[8][8] , \regs[8][7] , \regs[8][6] ,
         \regs[8][5] , \regs[8][4] , \regs[8][3] , \regs[8][2] , \regs[8][1] ,
         \regs[8][0] , \regs[7][15] , \regs[7][14] , \regs[7][13] ,
         \regs[7][12] , \regs[7][11] , \regs[7][10] , \regs[7][9] ,
         \regs[7][8] , \regs[7][7] , \regs[7][6] , \regs[7][5] , \regs[7][4] ,
         \regs[7][3] , \regs[7][2] , \regs[7][1] , \regs[7][0] , \regs[6][15] ,
         \regs[6][14] , \regs[6][13] , \regs[6][12] , \regs[6][11] ,
         \regs[6][10] , \regs[6][9] , \regs[6][8] , \regs[6][7] , \regs[6][6] ,
         \regs[6][5] , \regs[6][4] , \regs[6][3] , \regs[6][2] , \regs[6][1] ,
         \regs[6][0] , \regs[5][15] , \regs[5][14] , \regs[5][13] ,
         \regs[5][12] , \regs[5][11] , \regs[5][10] , \regs[5][9] ,
         \regs[5][8] , \regs[5][7] , \regs[5][6] , \regs[5][5] , \regs[5][4] ,
         \regs[5][3] , \regs[5][2] , \regs[5][1] , \regs[5][0] , \regs[4][15] ,
         \regs[4][14] , \regs[4][13] , \regs[4][12] , \regs[4][11] ,
         \regs[4][10] , \regs[4][9] , \regs[4][8] , \regs[4][7] , \regs[4][6] ,
         \regs[4][5] , \regs[4][4] , \regs[4][3] , \regs[4][2] , \regs[4][1] ,
         \regs[4][0] , \regs[3][15] , \regs[3][14] , \regs[3][13] ,
         \regs[3][12] , \regs[3][11] , \regs[3][10] , \regs[3][9] ,
         \regs[3][8] , \regs[3][7] , \regs[3][6] , \regs[3][5] , \regs[3][4] ,
         \regs[3][3] , \regs[3][2] , \regs[3][1] , \regs[3][0] , \regs[2][15] ,
         \regs[2][14] , \regs[2][13] , \regs[2][12] , \regs[2][11] ,
         \regs[2][10] , \regs[2][9] , \regs[2][8] , \regs[2][7] , \regs[2][6] ,
         \regs[2][5] , \regs[2][4] , \regs[2][3] , \regs[2][2] , \regs[2][1] ,
         \regs[2][0] , \regs[1][15] , \regs[1][14] , \regs[1][13] ,
         \regs[1][12] , \regs[1][11] , \regs[1][10] , \regs[1][9] ,
         \regs[1][8] , \regs[1][7] , \regs[1][6] , \regs[1][5] , \regs[1][4] ,
         \regs[1][3] , \regs[1][2] , \regs[1][1] , \regs[1][0] , n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n554, n769, n985, n993, n995, n999,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1017, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n986, n987, n988, n989,
         n990, n991, n992, n994, n996, n997, n998, n1000, n1016, n1018, n1035,
         n1053, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578;

  DFFSR \regs_reg[15][15]  ( .D(n257), .CLK(clk), .R(n599), .S(1'b1), .Q(
        \regs[15][15] ) );
  DFFSR \regs_reg[15][14]  ( .D(n258), .CLK(clk), .R(n599), .S(1'b1), .Q(
        \regs[15][14] ) );
  DFFSR \regs_reg[15][13]  ( .D(n259), .CLK(clk), .R(n599), .S(1'b1), .Q(
        \regs[15][13] ) );
  DFFSR \regs_reg[15][12]  ( .D(n260), .CLK(clk), .R(n599), .S(1'b1), .Q(
        \regs[15][12] ) );
  DFFSR \regs_reg[15][11]  ( .D(n261), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][11] ) );
  DFFSR \regs_reg[15][10]  ( .D(n262), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][10] ) );
  DFFSR \regs_reg[15][9]  ( .D(n263), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][9] ) );
  DFFSR \regs_reg[15][8]  ( .D(n264), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][8] ) );
  DFFSR \regs_reg[15][7]  ( .D(n265), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][7] ) );
  DFFSR \regs_reg[15][6]  ( .D(n266), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][6] ) );
  DFFSR \regs_reg[15][5]  ( .D(n267), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][5] ) );
  DFFSR \regs_reg[15][4]  ( .D(n268), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][4] ) );
  DFFSR \regs_reg[15][3]  ( .D(n269), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][3] ) );
  DFFSR \regs_reg[15][2]  ( .D(n270), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][2] ) );
  DFFSR \regs_reg[15][1]  ( .D(n271), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][1] ) );
  DFFSR \regs_reg[15][0]  ( .D(n272), .CLK(clk), .R(n598), .S(1'b1), .Q(
        \regs[15][0] ) );
  DFFSR \regs_reg[14][15]  ( .D(n273), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][15] ) );
  DFFSR \regs_reg[14][14]  ( .D(n274), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][14] ) );
  DFFSR \regs_reg[14][13]  ( .D(n275), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][13] ) );
  DFFSR \regs_reg[14][12]  ( .D(n276), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][12] ) );
  DFFSR \regs_reg[14][11]  ( .D(n277), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][11] ) );
  DFFSR \regs_reg[14][10]  ( .D(n278), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][10] ) );
  DFFSR \regs_reg[14][9]  ( .D(n279), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][9] ) );
  DFFSR \regs_reg[14][8]  ( .D(n280), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][8] ) );
  DFFSR \regs_reg[14][7]  ( .D(n281), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][7] ) );
  DFFSR \regs_reg[14][6]  ( .D(n282), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][6] ) );
  DFFSR \regs_reg[14][5]  ( .D(n283), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][5] ) );
  DFFSR \regs_reg[14][4]  ( .D(n284), .CLK(clk), .R(n597), .S(1'b1), .Q(
        \regs[14][4] ) );
  DFFSR \regs_reg[14][3]  ( .D(n285), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[14][3] ) );
  DFFSR \regs_reg[14][2]  ( .D(n286), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[14][2] ) );
  DFFSR \regs_reg[14][1]  ( .D(n287), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[14][1] ) );
  DFFSR \regs_reg[14][0]  ( .D(n288), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[14][0] ) );
  DFFSR \regs_reg[13][15]  ( .D(n289), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][15] ) );
  DFFSR \regs_reg[13][14]  ( .D(n290), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][14] ) );
  DFFSR \regs_reg[13][13]  ( .D(n291), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][13] ) );
  DFFSR \regs_reg[13][12]  ( .D(n292), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][12] ) );
  DFFSR \regs_reg[13][11]  ( .D(n293), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][11] ) );
  DFFSR \regs_reg[13][10]  ( .D(n294), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][10] ) );
  DFFSR \regs_reg[13][9]  ( .D(n295), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][9] ) );
  DFFSR \regs_reg[13][8]  ( .D(n296), .CLK(clk), .R(n596), .S(1'b1), .Q(
        \regs[13][8] ) );
  DFFSR \regs_reg[13][7]  ( .D(n297), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][7] ) );
  DFFSR \regs_reg[13][6]  ( .D(n298), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][6] ) );
  DFFSR \regs_reg[13][5]  ( .D(n299), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][5] ) );
  DFFSR \regs_reg[13][4]  ( .D(n300), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][4] ) );
  DFFSR \regs_reg[13][3]  ( .D(n301), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][3] ) );
  DFFSR \regs_reg[13][2]  ( .D(n302), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][2] ) );
  DFFSR \regs_reg[13][1]  ( .D(n303), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][1] ) );
  DFFSR \regs_reg[13][0]  ( .D(n304), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[13][0] ) );
  DFFSR \regs_reg[12][15]  ( .D(n305), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[12][15] ) );
  DFFSR \regs_reg[12][14]  ( .D(n306), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[12][14] ) );
  DFFSR \regs_reg[12][13]  ( .D(n307), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[12][13] ) );
  DFFSR \regs_reg[12][12]  ( .D(n308), .CLK(clk), .R(n595), .S(1'b1), .Q(
        \regs[12][12] ) );
  DFFSR \regs_reg[12][11]  ( .D(n309), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][11] ) );
  DFFSR \regs_reg[12][10]  ( .D(n310), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][10] ) );
  DFFSR \regs_reg[12][9]  ( .D(n311), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][9] ) );
  DFFSR \regs_reg[12][8]  ( .D(n312), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][8] ) );
  DFFSR \regs_reg[12][7]  ( .D(n313), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][7] ) );
  DFFSR \regs_reg[12][6]  ( .D(n314), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][6] ) );
  DFFSR \regs_reg[12][5]  ( .D(n315), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][5] ) );
  DFFSR \regs_reg[12][4]  ( .D(n316), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][4] ) );
  DFFSR \regs_reg[12][3]  ( .D(n317), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][3] ) );
  DFFSR \regs_reg[12][2]  ( .D(n318), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][2] ) );
  DFFSR \regs_reg[12][1]  ( .D(n319), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][1] ) );
  DFFSR \regs_reg[12][0]  ( .D(n320), .CLK(clk), .R(n594), .S(1'b1), .Q(
        \regs[12][0] ) );
  DFFSR \regs_reg[11][15]  ( .D(n1268), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][15] ) );
  DFFSR \regs_reg[11][14]  ( .D(n1267), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][14] ) );
  DFFSR \regs_reg[11][13]  ( .D(n1266), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][13] ) );
  DFFSR \regs_reg[11][12]  ( .D(n1265), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][12] ) );
  DFFSR \regs_reg[11][11]  ( .D(n1264), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][11] ) );
  DFFSR \regs_reg[11][10]  ( .D(n1263), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][10] ) );
  DFFSR \regs_reg[11][9]  ( .D(n1262), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][9] ) );
  DFFSR \regs_reg[11][8]  ( .D(n1261), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][8] ) );
  DFFSR \regs_reg[11][7]  ( .D(n1260), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][7] ) );
  DFFSR \regs_reg[11][6]  ( .D(n1259), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][6] ) );
  DFFSR \regs_reg[11][5]  ( .D(n1258), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][5] ) );
  DFFSR \regs_reg[11][4]  ( .D(n1257), .CLK(clk), .R(n593), .S(1'b1), .Q(
        \regs[11][4] ) );
  DFFSR \regs_reg[11][3]  ( .D(n1256), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[11][3] ) );
  DFFSR \regs_reg[11][2]  ( .D(n1255), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[11][2] ) );
  DFFSR \regs_reg[11][1]  ( .D(n1254), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[11][1] ) );
  DFFSR \regs_reg[11][0]  ( .D(n1253), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[11][0] ) );
  DFFSR \regs_reg[10][15]  ( .D(n1252), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][15] ) );
  DFFSR \regs_reg[10][14]  ( .D(n1251), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][14] ) );
  DFFSR \regs_reg[10][13]  ( .D(n1250), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][13] ) );
  DFFSR \regs_reg[10][12]  ( .D(n1249), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][12] ) );
  DFFSR \regs_reg[10][11]  ( .D(n1248), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][11] ) );
  DFFSR \regs_reg[10][10]  ( .D(n1247), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][10] ) );
  DFFSR \regs_reg[10][9]  ( .D(n1246), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][9] ) );
  DFFSR \regs_reg[10][8]  ( .D(n1245), .CLK(clk), .R(n592), .S(1'b1), .Q(
        \regs[10][8] ) );
  DFFSR \regs_reg[10][7]  ( .D(n1244), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][7] ) );
  DFFSR \regs_reg[10][6]  ( .D(n1243), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][6] ) );
  DFFSR \regs_reg[10][5]  ( .D(n1242), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][5] ) );
  DFFSR \regs_reg[10][4]  ( .D(n1241), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][4] ) );
  DFFSR \regs_reg[10][3]  ( .D(n1240), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][3] ) );
  DFFSR \regs_reg[10][2]  ( .D(n1239), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][2] ) );
  DFFSR \regs_reg[10][1]  ( .D(n1238), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][1] ) );
  DFFSR \regs_reg[10][0]  ( .D(n1237), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[10][0] ) );
  DFFSR \regs_reg[9][15]  ( .D(n1236), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[9][15] ) );
  DFFSR \regs_reg[9][14]  ( .D(n1235), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[9][14] ) );
  DFFSR \regs_reg[9][13]  ( .D(n1234), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[9][13] ) );
  DFFSR \regs_reg[9][12]  ( .D(n1233), .CLK(clk), .R(n591), .S(1'b1), .Q(
        \regs[9][12] ) );
  DFFSR \regs_reg[9][11]  ( .D(n1232), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][11] ) );
  DFFSR \regs_reg[9][10]  ( .D(n1231), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][10] ) );
  DFFSR \regs_reg[9][9]  ( .D(n1230), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][9] ) );
  DFFSR \regs_reg[9][8]  ( .D(n1229), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][8] ) );
  DFFSR \regs_reg[9][7]  ( .D(n1228), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][7] ) );
  DFFSR \regs_reg[9][6]  ( .D(n1227), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][6] ) );
  DFFSR \regs_reg[9][5]  ( .D(n1226), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][5] ) );
  DFFSR \regs_reg[9][4]  ( .D(n1225), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][4] ) );
  DFFSR \regs_reg[9][3]  ( .D(n1224), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][3] ) );
  DFFSR \regs_reg[9][2]  ( .D(n1223), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][2] ) );
  DFFSR \regs_reg[9][1]  ( .D(n1222), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][1] ) );
  DFFSR \regs_reg[9][0]  ( .D(n1221), .CLK(clk), .R(n590), .S(1'b1), .Q(
        \regs[9][0] ) );
  DFFSR \regs_reg[8][15]  ( .D(n1220), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][15] ) );
  DFFSR \regs_reg[8][14]  ( .D(n1219), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][14] ) );
  DFFSR \regs_reg[8][13]  ( .D(n1218), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][13] ) );
  DFFSR \regs_reg[8][12]  ( .D(n1217), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][12] ) );
  DFFSR \regs_reg[8][11]  ( .D(n1216), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][11] ) );
  DFFSR \regs_reg[8][10]  ( .D(n1215), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][10] ) );
  DFFSR \regs_reg[8][9]  ( .D(n1214), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][9] ) );
  DFFSR \regs_reg[8][8]  ( .D(n1213), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][8] ) );
  DFFSR \regs_reg[8][7]  ( .D(n1212), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][7] ) );
  DFFSR \regs_reg[8][6]  ( .D(n1211), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][6] ) );
  DFFSR \regs_reg[8][5]  ( .D(n1210), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][5] ) );
  DFFSR \regs_reg[8][4]  ( .D(n1209), .CLK(clk), .R(n589), .S(1'b1), .Q(
        \regs[8][4] ) );
  DFFSR \regs_reg[8][3]  ( .D(n1208), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[8][3] ) );
  DFFSR \regs_reg[8][2]  ( .D(n1207), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[8][2] ) );
  DFFSR \regs_reg[8][1]  ( .D(n1206), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[8][1] ) );
  DFFSR \regs_reg[8][0]  ( .D(n1205), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[8][0] ) );
  DFFSR \regs_reg[7][15]  ( .D(n1204), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][15] ) );
  DFFSR \regs_reg[7][14]  ( .D(n1203), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][14] ) );
  DFFSR \regs_reg[7][13]  ( .D(n1202), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][13] ) );
  DFFSR \regs_reg[7][12]  ( .D(n1201), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][12] ) );
  DFFSR \regs_reg[7][11]  ( .D(n1200), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][11] ) );
  DFFSR \regs_reg[7][10]  ( .D(n1199), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][10] ) );
  DFFSR \regs_reg[7][9]  ( .D(n1198), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][9] ) );
  DFFSR \regs_reg[7][8]  ( .D(n1197), .CLK(clk), .R(n588), .S(1'b1), .Q(
        \regs[7][8] ) );
  DFFSR \regs_reg[7][7]  ( .D(n1196), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][7] ) );
  DFFSR \regs_reg[7][6]  ( .D(n1195), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][6] ) );
  DFFSR \regs_reg[7][5]  ( .D(n1194), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][5] ) );
  DFFSR \regs_reg[7][4]  ( .D(n1193), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][4] ) );
  DFFSR \regs_reg[7][3]  ( .D(n1192), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][3] ) );
  DFFSR \regs_reg[7][2]  ( .D(n1191), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][2] ) );
  DFFSR \regs_reg[7][1]  ( .D(n1190), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][1] ) );
  DFFSR \regs_reg[7][0]  ( .D(n1189), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[7][0] ) );
  DFFSR \regs_reg[6][15]  ( .D(n1188), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[6][15] ) );
  DFFSR \regs_reg[6][14]  ( .D(n1187), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[6][14] ) );
  DFFSR \regs_reg[6][13]  ( .D(n1186), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[6][13] ) );
  DFFSR \regs_reg[6][12]  ( .D(n1185), .CLK(clk), .R(n587), .S(1'b1), .Q(
        \regs[6][12] ) );
  DFFSR \regs_reg[6][11]  ( .D(n1184), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][11] ) );
  DFFSR \regs_reg[6][10]  ( .D(n1183), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][10] ) );
  DFFSR \regs_reg[6][9]  ( .D(n1182), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][9] ) );
  DFFSR \regs_reg[6][8]  ( .D(n1181), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][8] ) );
  DFFSR \regs_reg[6][7]  ( .D(n1180), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][7] ) );
  DFFSR \regs_reg[6][6]  ( .D(n1179), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][6] ) );
  DFFSR \regs_reg[6][5]  ( .D(n1178), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][5] ) );
  DFFSR \regs_reg[6][4]  ( .D(n1177), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][4] ) );
  DFFSR \regs_reg[6][3]  ( .D(n1176), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][3] ) );
  DFFSR \regs_reg[6][2]  ( .D(n1175), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][2] ) );
  DFFSR \regs_reg[6][1]  ( .D(n1174), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][1] ) );
  DFFSR \regs_reg[6][0]  ( .D(n1173), .CLK(clk), .R(n586), .S(1'b1), .Q(
        \regs[6][0] ) );
  DFFSR \regs_reg[5][15]  ( .D(n1172), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][15] ) );
  DFFSR \regs_reg[5][14]  ( .D(n1171), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][14] ) );
  DFFSR \regs_reg[5][13]  ( .D(n1170), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][13] ) );
  DFFSR \regs_reg[5][12]  ( .D(n1169), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][12] ) );
  DFFSR \regs_reg[5][11]  ( .D(n1168), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][11] ) );
  DFFSR \regs_reg[5][10]  ( .D(n1167), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][10] ) );
  DFFSR \regs_reg[5][9]  ( .D(n1166), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][9] ) );
  DFFSR \regs_reg[5][8]  ( .D(n1165), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][8] ) );
  DFFSR \regs_reg[5][7]  ( .D(n1164), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][7] ) );
  DFFSR \regs_reg[5][6]  ( .D(n1163), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][6] ) );
  DFFSR \regs_reg[5][5]  ( .D(n1162), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][5] ) );
  DFFSR \regs_reg[5][4]  ( .D(n1161), .CLK(clk), .R(n585), .S(1'b1), .Q(
        \regs[5][4] ) );
  DFFSR \regs_reg[5][3]  ( .D(n1160), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[5][3] ) );
  DFFSR \regs_reg[5][2]  ( .D(n1159), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[5][2] ) );
  DFFSR \regs_reg[5][1]  ( .D(n1158), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[5][1] ) );
  DFFSR \regs_reg[5][0]  ( .D(n1157), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[5][0] ) );
  DFFSR \regs_reg[4][15]  ( .D(n1156), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][15] ) );
  DFFSR \regs_reg[4][14]  ( .D(n1155), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][14] ) );
  DFFSR \regs_reg[4][13]  ( .D(n1154), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][13] ) );
  DFFSR \regs_reg[4][12]  ( .D(n1153), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][12] ) );
  DFFSR \regs_reg[4][11]  ( .D(n1152), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][11] ) );
  DFFSR \regs_reg[4][10]  ( .D(n1151), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][10] ) );
  DFFSR \regs_reg[4][9]  ( .D(n1150), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][9] ) );
  DFFSR \regs_reg[4][8]  ( .D(n1149), .CLK(clk), .R(n584), .S(1'b1), .Q(
        \regs[4][8] ) );
  DFFSR \regs_reg[4][7]  ( .D(n1148), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][7] ) );
  DFFSR \regs_reg[4][6]  ( .D(n1147), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][6] ) );
  DFFSR \regs_reg[4][5]  ( .D(n1146), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][5] ) );
  DFFSR \regs_reg[4][4]  ( .D(n1145), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][4] ) );
  DFFSR \regs_reg[4][3]  ( .D(n1144), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][3] ) );
  DFFSR \regs_reg[4][2]  ( .D(n1143), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][2] ) );
  DFFSR \regs_reg[4][1]  ( .D(n1142), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][1] ) );
  DFFSR \regs_reg[4][0]  ( .D(n1141), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[4][0] ) );
  DFFSR \regs_reg[3][15]  ( .D(n449), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[3][15] ) );
  DFFSR \regs_reg[3][14]  ( .D(n450), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[3][14] ) );
  DFFSR \regs_reg[3][13]  ( .D(n451), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[3][13] ) );
  DFFSR \regs_reg[3][12]  ( .D(n452), .CLK(clk), .R(n583), .S(1'b1), .Q(
        \regs[3][12] ) );
  DFFSR \regs_reg[3][11]  ( .D(n453), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][11] ) );
  DFFSR \regs_reg[3][10]  ( .D(n454), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][10] ) );
  DFFSR \regs_reg[3][9]  ( .D(n455), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][9] ) );
  DFFSR \regs_reg[3][8]  ( .D(n456), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][8] ) );
  DFFSR \regs_reg[3][7]  ( .D(n457), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][7] ) );
  DFFSR \regs_reg[3][6]  ( .D(n458), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][6] ) );
  DFFSR \regs_reg[3][5]  ( .D(n459), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][5] ) );
  DFFSR \regs_reg[3][4]  ( .D(n460), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][4] ) );
  DFFSR \regs_reg[3][3]  ( .D(n461), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][3] ) );
  DFFSR \regs_reg[3][2]  ( .D(n462), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][2] ) );
  DFFSR \regs_reg[3][1]  ( .D(n463), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][1] ) );
  DFFSR \regs_reg[3][0]  ( .D(n464), .CLK(clk), .R(n582), .S(1'b1), .Q(
        \regs[3][0] ) );
  DFFSR \regs_reg[2][15]  ( .D(n465), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][15] ) );
  DFFSR \regs_reg[2][14]  ( .D(n466), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][14] ) );
  DFFSR \regs_reg[2][13]  ( .D(n467), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][13] ) );
  DFFSR \regs_reg[2][12]  ( .D(n468), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][12] ) );
  DFFSR \regs_reg[2][11]  ( .D(n469), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][11] ) );
  DFFSR \regs_reg[2][10]  ( .D(n470), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][10] ) );
  DFFSR \regs_reg[2][9]  ( .D(n471), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][9] ) );
  DFFSR \regs_reg[2][8]  ( .D(n472), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][8] ) );
  DFFSR \regs_reg[2][7]  ( .D(n473), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][7] ) );
  DFFSR \regs_reg[2][6]  ( .D(n474), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][6] ) );
  DFFSR \regs_reg[2][5]  ( .D(n475), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][5] ) );
  DFFSR \regs_reg[2][4]  ( .D(n476), .CLK(clk), .R(n581), .S(1'b1), .Q(
        \regs[2][4] ) );
  DFFSR \regs_reg[2][3]  ( .D(n477), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[2][3] ) );
  DFFSR \regs_reg[2][2]  ( .D(n478), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[2][2] ) );
  DFFSR \regs_reg[2][1]  ( .D(n479), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[2][1] ) );
  DFFSR \regs_reg[2][0]  ( .D(n480), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[2][0] ) );
  DFFSR \regs_reg[1][15]  ( .D(n481), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][15] ) );
  DFFSR \regs_reg[1][14]  ( .D(n482), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][14] ) );
  DFFSR \regs_reg[1][13]  ( .D(n483), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][13] ) );
  DFFSR \regs_reg[1][12]  ( .D(n484), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][12] ) );
  DFFSR \regs_reg[1][11]  ( .D(n485), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][11] ) );
  DFFSR \regs_reg[1][10]  ( .D(n486), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][10] ) );
  DFFSR \regs_reg[1][9]  ( .D(n487), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][9] ) );
  DFFSR \regs_reg[1][8]  ( .D(n488), .CLK(clk), .R(n580), .S(1'b1), .Q(
        \regs[1][8] ) );
  DFFSR \regs_reg[1][7]  ( .D(n489), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][7] ) );
  DFFSR \regs_reg[1][6]  ( .D(n490), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][6] ) );
  DFFSR \regs_reg[1][5]  ( .D(n491), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][5] ) );
  DFFSR \regs_reg[1][4]  ( .D(n492), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][4] ) );
  DFFSR \regs_reg[1][3]  ( .D(n493), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][3] ) );
  DFFSR \regs_reg[1][2]  ( .D(n494), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][2] ) );
  DFFSR \regs_reg[1][1]  ( .D(n495), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][1] ) );
  DFFSR \regs_reg[1][0]  ( .D(n496), .CLK(clk), .R(n579), .S(1'b1), .Q(
        \regs[1][0] ) );
  DFFSR \regs_reg[0][15]  ( .D(n497), .CLK(clk), .R(n579), .S(1'b1), .Q(
        outreg_data[15]) );
  DFFSR \regs_reg[0][14]  ( .D(n498), .CLK(clk), .R(n579), .S(1'b1), .Q(
        outreg_data[14]) );
  DFFSR \regs_reg[0][13]  ( .D(n499), .CLK(clk), .R(n579), .S(1'b1), .Q(
        outreg_data[13]) );
  DFFSR \regs_reg[0][12]  ( .D(n500), .CLK(clk), .R(n579), .S(1'b1), .Q(
        outreg_data[12]) );
  DFFSR \regs_reg[0][11]  ( .D(n501), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[11]) );
  DFFSR \regs_reg[0][10]  ( .D(n502), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[10]) );
  DFFSR \regs_reg[0][9]  ( .D(n503), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[9]) );
  DFFSR \regs_reg[0][8]  ( .D(n504), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[8]) );
  DFFSR \regs_reg[0][7]  ( .D(n505), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[7]) );
  DFFSR \regs_reg[0][6]  ( .D(n506), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[6]) );
  DFFSR \regs_reg[0][5]  ( .D(n507), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[5]) );
  DFFSR \regs_reg[0][4]  ( .D(n508), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[4]) );
  DFFSR \regs_reg[0][3]  ( .D(n509), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[3]) );
  DFFSR \regs_reg[0][2]  ( .D(n510), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[2]) );
  DFFSR \regs_reg[0][1]  ( .D(n511), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[1]) );
  DFFSR \regs_reg[0][0]  ( .D(n512), .CLK(clk), .R(n578), .S(1'b1), .Q(
        outreg_data[0]) );
  AND2X2 U310 ( .A(n1051), .B(n1578), .Y(n993) );
  AND2X2 U311 ( .A(n1051), .B(w_sel[0]), .Y(n995) );
  AND2X2 U312 ( .A(w_sel[3]), .B(w_en), .Y(n1051) );
  INVX2 U315 ( .A(n1068), .Y(n257) );
  INVX2 U316 ( .A(n1067), .Y(n258) );
  INVX2 U317 ( .A(n1066), .Y(n259) );
  INVX2 U318 ( .A(n1065), .Y(n260) );
  INVX2 U319 ( .A(n1064), .Y(n261) );
  INVX2 U320 ( .A(n1063), .Y(n262) );
  INVX2 U321 ( .A(n1062), .Y(n263) );
  INVX2 U322 ( .A(n1061), .Y(n264) );
  INVX2 U323 ( .A(n1060), .Y(n265) );
  INVX2 U324 ( .A(n1059), .Y(n266) );
  INVX2 U325 ( .A(n1058), .Y(n267) );
  INVX2 U326 ( .A(n1057), .Y(n268) );
  INVX2 U327 ( .A(n1056), .Y(n269) );
  INVX2 U328 ( .A(n1055), .Y(n270) );
  INVX2 U329 ( .A(n1054), .Y(n271) );
  INVX2 U330 ( .A(n1052), .Y(n272) );
  INVX2 U331 ( .A(n1050), .Y(n273) );
  INVX2 U332 ( .A(n1049), .Y(n274) );
  INVX2 U333 ( .A(n1048), .Y(n275) );
  INVX2 U334 ( .A(n1047), .Y(n276) );
  INVX2 U335 ( .A(n1046), .Y(n277) );
  INVX2 U336 ( .A(n1045), .Y(n278) );
  INVX2 U337 ( .A(n1044), .Y(n279) );
  INVX2 U338 ( .A(n1043), .Y(n280) );
  INVX2 U339 ( .A(n1042), .Y(n281) );
  INVX2 U340 ( .A(n1041), .Y(n282) );
  INVX2 U341 ( .A(n1040), .Y(n283) );
  INVX2 U342 ( .A(n1039), .Y(n284) );
  INVX2 U343 ( .A(n1038), .Y(n285) );
  INVX2 U344 ( .A(n1037), .Y(n286) );
  INVX2 U345 ( .A(n1036), .Y(n287) );
  INVX2 U346 ( .A(n1034), .Y(n288) );
  INVX2 U347 ( .A(n1033), .Y(n289) );
  INVX2 U348 ( .A(n1032), .Y(n290) );
  INVX2 U349 ( .A(n1031), .Y(n291) );
  INVX2 U350 ( .A(n1030), .Y(n292) );
  INVX2 U351 ( .A(n1029), .Y(n293) );
  INVX2 U352 ( .A(n1028), .Y(n294) );
  INVX2 U353 ( .A(n1027), .Y(n295) );
  INVX2 U354 ( .A(n1026), .Y(n296) );
  INVX2 U355 ( .A(n1025), .Y(n297) );
  INVX2 U356 ( .A(n1024), .Y(n298) );
  INVX2 U357 ( .A(n1023), .Y(n299) );
  INVX2 U358 ( .A(n1022), .Y(n300) );
  INVX2 U359 ( .A(n1021), .Y(n301) );
  INVX2 U360 ( .A(n1020), .Y(n302) );
  INVX2 U361 ( .A(n1019), .Y(n303) );
  INVX2 U362 ( .A(n1017), .Y(n304) );
  INVX2 U363 ( .A(n1015), .Y(n305) );
  INVX2 U364 ( .A(n1014), .Y(n306) );
  INVX2 U365 ( .A(n1013), .Y(n307) );
  INVX2 U366 ( .A(n1012), .Y(n308) );
  INVX2 U367 ( .A(n1011), .Y(n309) );
  INVX2 U368 ( .A(n1010), .Y(n310) );
  INVX2 U369 ( .A(n1009), .Y(n311) );
  INVX2 U370 ( .A(n1008), .Y(n312) );
  INVX2 U371 ( .A(n1007), .Y(n313) );
  INVX2 U372 ( .A(n1006), .Y(n314) );
  INVX2 U373 ( .A(n1005), .Y(n315) );
  INVX2 U374 ( .A(n1004), .Y(n316) );
  INVX2 U375 ( .A(n1003), .Y(n317) );
  INVX2 U376 ( .A(n1002), .Y(n318) );
  INVX2 U377 ( .A(n1001), .Y(n319) );
  INVX2 U378 ( .A(n999), .Y(n320) );
  INVX2 U612 ( .A(w_en), .Y(n554) );
  NOR2X1 U813 ( .A(n647), .B(n413), .Y(n769) );
  NOR2X1 U1019 ( .A(n1071), .B(n344), .Y(n985) );
  AOI22X1 U1120 ( .A(w_data[0]), .B(n526), .C(n569), .D(\regs[12][0] ), .Y(
        n999) );
  AOI22X1 U1121 ( .A(w_data[1]), .B(n526), .C(n569), .D(\regs[12][1] ), .Y(
        n1001) );
  AOI22X1 U1122 ( .A(w_data[2]), .B(n526), .C(n569), .D(\regs[12][2] ), .Y(
        n1002) );
  AOI22X1 U1123 ( .A(w_data[3]), .B(n526), .C(n569), .D(\regs[12][3] ), .Y(
        n1003) );
  AOI22X1 U1124 ( .A(w_data[4]), .B(n526), .C(n569), .D(\regs[12][4] ), .Y(
        n1004) );
  AOI22X1 U1125 ( .A(w_data[5]), .B(n526), .C(n569), .D(\regs[12][5] ), .Y(
        n1005) );
  AOI22X1 U1126 ( .A(w_data[6]), .B(n526), .C(n569), .D(\regs[12][6] ), .Y(
        n1006) );
  AOI22X1 U1127 ( .A(w_data[7]), .B(n526), .C(n569), .D(\regs[12][7] ), .Y(
        n1007) );
  AOI22X1 U1128 ( .A(w_data[8]), .B(n526), .C(n569), .D(\regs[12][8] ), .Y(
        n1008) );
  AOI22X1 U1129 ( .A(w_data[9]), .B(n526), .C(n569), .D(\regs[12][9] ), .Y(
        n1009) );
  AOI22X1 U1130 ( .A(w_data[10]), .B(n526), .C(n569), .D(\regs[12][10] ), .Y(
        n1010) );
  AOI22X1 U1131 ( .A(w_data[11]), .B(n526), .C(n569), .D(\regs[12][11] ), .Y(
        n1011) );
  AOI22X1 U1132 ( .A(w_data[12]), .B(n526), .C(n569), .D(\regs[12][12] ), .Y(
        n1012) );
  AOI22X1 U1133 ( .A(w_data[13]), .B(n526), .C(n569), .D(\regs[12][13] ), .Y(
        n1013) );
  AOI22X1 U1134 ( .A(w_data[14]), .B(n526), .C(n569), .D(\regs[12][14] ), .Y(
        n1014) );
  AOI22X1 U1135 ( .A(w_data[15]), .B(n526), .C(n569), .D(\regs[12][15] ), .Y(
        n1015) );
  AOI22X1 U1137 ( .A(w_data[0]), .B(n527), .C(n568), .D(\regs[13][0] ), .Y(
        n1017) );
  AOI22X1 U1138 ( .A(w_data[1]), .B(n527), .C(n568), .D(\regs[13][1] ), .Y(
        n1019) );
  AOI22X1 U1139 ( .A(w_data[2]), .B(n527), .C(n568), .D(\regs[13][2] ), .Y(
        n1020) );
  AOI22X1 U1140 ( .A(w_data[3]), .B(n527), .C(n568), .D(\regs[13][3] ), .Y(
        n1021) );
  AOI22X1 U1141 ( .A(w_data[4]), .B(n527), .C(n568), .D(\regs[13][4] ), .Y(
        n1022) );
  AOI22X1 U1142 ( .A(w_data[5]), .B(n527), .C(n568), .D(\regs[13][5] ), .Y(
        n1023) );
  AOI22X1 U1143 ( .A(w_data[6]), .B(n527), .C(n568), .D(\regs[13][6] ), .Y(
        n1024) );
  AOI22X1 U1144 ( .A(w_data[7]), .B(n527), .C(n568), .D(\regs[13][7] ), .Y(
        n1025) );
  AOI22X1 U1145 ( .A(w_data[8]), .B(n527), .C(n568), .D(\regs[13][8] ), .Y(
        n1026) );
  AOI22X1 U1146 ( .A(w_data[9]), .B(n527), .C(n568), .D(\regs[13][9] ), .Y(
        n1027) );
  AOI22X1 U1147 ( .A(w_data[10]), .B(n527), .C(n568), .D(\regs[13][10] ), .Y(
        n1028) );
  AOI22X1 U1148 ( .A(w_data[11]), .B(n527), .C(n568), .D(\regs[13][11] ), .Y(
        n1029) );
  AOI22X1 U1149 ( .A(w_data[12]), .B(n527), .C(n568), .D(\regs[13][12] ), .Y(
        n1030) );
  AOI22X1 U1150 ( .A(w_data[13]), .B(n527), .C(n568), .D(\regs[13][13] ), .Y(
        n1031) );
  AOI22X1 U1151 ( .A(w_data[14]), .B(n527), .C(n568), .D(\regs[13][14] ), .Y(
        n1032) );
  AOI22X1 U1152 ( .A(w_data[15]), .B(n527), .C(n568), .D(\regs[13][15] ), .Y(
        n1033) );
  AOI22X1 U1154 ( .A(w_data[0]), .B(n528), .C(n567), .D(\regs[14][0] ), .Y(
        n1034) );
  AOI22X1 U1155 ( .A(w_data[1]), .B(n528), .C(n567), .D(\regs[14][1] ), .Y(
        n1036) );
  AOI22X1 U1156 ( .A(w_data[2]), .B(n528), .C(n567), .D(\regs[14][2] ), .Y(
        n1037) );
  AOI22X1 U1157 ( .A(w_data[3]), .B(n528), .C(n567), .D(\regs[14][3] ), .Y(
        n1038) );
  AOI22X1 U1158 ( .A(w_data[4]), .B(n528), .C(n567), .D(\regs[14][4] ), .Y(
        n1039) );
  AOI22X1 U1159 ( .A(w_data[5]), .B(n528), .C(n567), .D(\regs[14][5] ), .Y(
        n1040) );
  AOI22X1 U1160 ( .A(w_data[6]), .B(n528), .C(n567), .D(\regs[14][6] ), .Y(
        n1041) );
  AOI22X1 U1161 ( .A(w_data[7]), .B(n528), .C(n567), .D(\regs[14][7] ), .Y(
        n1042) );
  AOI22X1 U1162 ( .A(w_data[8]), .B(n528), .C(n567), .D(\regs[14][8] ), .Y(
        n1043) );
  AOI22X1 U1163 ( .A(w_data[9]), .B(n528), .C(n567), .D(\regs[14][9] ), .Y(
        n1044) );
  AOI22X1 U1164 ( .A(w_data[10]), .B(n528), .C(n567), .D(\regs[14][10] ), .Y(
        n1045) );
  AOI22X1 U1165 ( .A(w_data[11]), .B(n528), .C(n567), .D(\regs[14][11] ), .Y(
        n1046) );
  AOI22X1 U1166 ( .A(w_data[12]), .B(n528), .C(n567), .D(\regs[14][12] ), .Y(
        n1047) );
  AOI22X1 U1167 ( .A(w_data[13]), .B(n528), .C(n567), .D(\regs[14][13] ), .Y(
        n1048) );
  AOI22X1 U1168 ( .A(w_data[14]), .B(n528), .C(n567), .D(\regs[14][14] ), .Y(
        n1049) );
  AOI22X1 U1169 ( .A(w_data[15]), .B(n528), .C(n567), .D(\regs[14][15] ), .Y(
        n1050) );
  AOI22X1 U1171 ( .A(w_data[0]), .B(n529), .C(n566), .D(\regs[15][0] ), .Y(
        n1052) );
  AOI22X1 U1172 ( .A(w_data[1]), .B(n529), .C(n566), .D(\regs[15][1] ), .Y(
        n1054) );
  AOI22X1 U1173 ( .A(w_data[2]), .B(n529), .C(n566), .D(\regs[15][2] ), .Y(
        n1055) );
  AOI22X1 U1174 ( .A(w_data[3]), .B(n529), .C(n566), .D(\regs[15][3] ), .Y(
        n1056) );
  AOI22X1 U1175 ( .A(w_data[4]), .B(n529), .C(n566), .D(\regs[15][4] ), .Y(
        n1057) );
  AOI22X1 U1176 ( .A(w_data[5]), .B(n529), .C(n566), .D(\regs[15][5] ), .Y(
        n1058) );
  AOI22X1 U1177 ( .A(w_data[6]), .B(n529), .C(n566), .D(\regs[15][6] ), .Y(
        n1059) );
  AOI22X1 U1178 ( .A(w_data[7]), .B(n529), .C(n566), .D(\regs[15][7] ), .Y(
        n1060) );
  AOI22X1 U1179 ( .A(w_data[8]), .B(n529), .C(n566), .D(\regs[15][8] ), .Y(
        n1061) );
  AOI22X1 U1180 ( .A(w_data[9]), .B(n529), .C(n566), .D(\regs[15][9] ), .Y(
        n1062) );
  AOI22X1 U1181 ( .A(w_data[10]), .B(n529), .C(n566), .D(\regs[15][10] ), .Y(
        n1063) );
  AOI22X1 U1182 ( .A(w_data[11]), .B(n529), .C(n566), .D(\regs[15][11] ), .Y(
        n1064) );
  AOI22X1 U1183 ( .A(w_data[12]), .B(n529), .C(n566), .D(\regs[15][12] ), .Y(
        n1065) );
  AOI22X1 U1184 ( .A(w_data[13]), .B(n529), .C(n566), .D(\regs[15][13] ), .Y(
        n1066) );
  AOI22X1 U1185 ( .A(w_data[14]), .B(n529), .C(n566), .D(\regs[15][14] ), .Y(
        n1067) );
  AOI22X1 U1186 ( .A(w_data[15]), .B(n529), .C(n566), .D(\regs[15][15] ), .Y(
        n1068) );
  NOR2X1 U1300 ( .A(n554), .B(w_sel[3]), .Y(n1140) );
  NAND2X1 U258 ( .A(n325), .B(n519), .Y(n321) );
  OR2X2 U259 ( .A(n1475), .B(r1_sel[0]), .Y(n1087) );
  BUFX4 U260 ( .A(n996), .Y(n322) );
  INVX2 U261 ( .A(r2_sel[2]), .Y(n345) );
  INVX1 U262 ( .A(n789), .Y(n323) );
  INVX2 U263 ( .A(n533), .Y(n324) );
  INVX2 U264 ( .A(n324), .Y(n325) );
  INVX2 U265 ( .A(w_data[11]), .Y(n326) );
  INVX2 U266 ( .A(r2_sel[2]), .Y(n351) );
  INVX1 U267 ( .A(w_data[8]), .Y(n327) );
  INVX2 U268 ( .A(w_data[6]), .Y(n328) );
  INVX2 U269 ( .A(w_data[5]), .Y(n329) );
  INVX1 U270 ( .A(w_data[12]), .Y(n330) );
  INVX1 U271 ( .A(w_data[10]), .Y(n334) );
  INVX1 U272 ( .A(w_data[15]), .Y(n335) );
  INVX2 U273 ( .A(w_data[9]), .Y(n331) );
  INVX1 U274 ( .A(w_data[14]), .Y(n336) );
  INVX1 U275 ( .A(n323), .Y(n431) );
  INVX2 U276 ( .A(w_data[11]), .Y(n332) );
  INVX1 U277 ( .A(n925), .Y(n333) );
  AND2X1 U278 ( .A(n1140), .B(n1578), .Y(n337) );
  AND2X1 U279 ( .A(n1140), .B(w_sel[0]), .Y(n338) );
  INVX4 U280 ( .A(n893), .Y(n430) );
  INVX4 U281 ( .A(n869), .Y(n410) );
  INVX2 U282 ( .A(r1_sel[0]), .Y(n391) );
  INVX1 U283 ( .A(n333), .Y(n347) );
  INVX2 U284 ( .A(n438), .Y(n339) );
  INVX4 U285 ( .A(n821), .Y(n438) );
  INVX2 U286 ( .A(r2_sel[1]), .Y(n821) );
  INVX4 U287 ( .A(n1422), .Y(n1560) );
  INVX4 U288 ( .A(n564), .Y(n1335) );
  INVX2 U289 ( .A(n410), .Y(n340) );
  INVX1 U290 ( .A(n775), .Y(n341) );
  INVX1 U291 ( .A(n775), .Y(n422) );
  INVX1 U292 ( .A(n396), .Y(n342) );
  INVX2 U293 ( .A(n396), .Y(n796) );
  INVX1 U294 ( .A(r1_sel[2]), .Y(n343) );
  INVX2 U295 ( .A(n343), .Y(n344) );
  INVX1 U296 ( .A(n345), .Y(n346) );
  INVX1 U297 ( .A(n423), .Y(n348) );
  INVX2 U298 ( .A(n892), .Y(n349) );
  INVX1 U299 ( .A(r2_sel[2]), .Y(n395) );
  OR2X1 U300 ( .A(n1069), .B(n1053), .Y(r2_data[15]) );
  NAND2X1 U301 ( .A(n1375), .B(r1_sel[1]), .Y(n350) );
  INVX2 U302 ( .A(n350), .Y(n417) );
  OR2X1 U303 ( .A(n831), .B(n832), .Y(r2_data[8]) );
  INVX4 U304 ( .A(n988), .Y(n425) );
  BUFX2 U305 ( .A(n514), .Y(n352) );
  INVX1 U306 ( .A(n989), .Y(n353) );
  INVX1 U307 ( .A(n513), .Y(n354) );
  INVX1 U308 ( .A(n354), .Y(n355) );
  INVX1 U309 ( .A(n342), .Y(n356) );
  INVX1 U313 ( .A(n796), .Y(n401) );
  INVX2 U314 ( .A(n551), .Y(n357) );
  AND2X2 U379 ( .A(n752), .B(n751), .Y(n362) );
  INVX4 U380 ( .A(n428), .Y(n358) );
  INVX2 U381 ( .A(n353), .Y(n429) );
  INVX2 U382 ( .A(n989), .Y(n428) );
  INVX4 U383 ( .A(n991), .Y(n550) );
  INVX2 U384 ( .A(n600), .Y(n603) );
  INVX2 U385 ( .A(n603), .Y(n372) );
  INVX2 U386 ( .A(n969), .Y(n370) );
  INVX4 U387 ( .A(n605), .Y(n969) );
  INVX2 U388 ( .A(n965), .Y(n371) );
  INVX2 U389 ( .A(n607), .Y(n965) );
  INVX2 U390 ( .A(n967), .Y(n369) );
  INVX2 U391 ( .A(n609), .Y(n967) );
  INVX2 U392 ( .A(\regs[5][10] ), .Y(n1444) );
  AND2X2 U393 ( .A(w_sel[1]), .B(w_sel[2]), .Y(n359) );
  AND2X2 U394 ( .A(w_sel[2]), .B(n613), .Y(n360) );
  AND2X2 U395 ( .A(n1438), .B(n1375), .Y(n361) );
  AND2X2 U396 ( .A(n993), .B(n359), .Y(n528) );
  INVX2 U397 ( .A(n868), .Y(n432) );
  AND2X1 U398 ( .A(n1427), .B(n1426), .Y(n363) );
  AND2X1 U399 ( .A(n1314), .B(n1313), .Y(n364) );
  AND2X2 U400 ( .A(n1140), .B(n618), .Y(n365) );
  AND2X2 U401 ( .A(n536), .B(n519), .Y(n366) );
  INVX8 U402 ( .A(w_data[1]), .Y(n645) );
  INVX2 U403 ( .A(w_data[4]), .Y(n367) );
  MUX2X1 U404 ( .B(n814), .A(n824), .S(n434), .Y(n1197) );
  MUX2X1 U405 ( .B(n814), .A(n825), .S(n437), .Y(n1181) );
  MUX2X1 U406 ( .B(n814), .A(n810), .S(n368), .Y(n1165) );
  MUX2X1 U407 ( .B(n814), .A(n811), .S(n435), .Y(n1149) );
  MUX2X1 U408 ( .B(n814), .A(n813), .S(n369), .Y(n456) );
  MUX2X1 U409 ( .B(n814), .A(n812), .S(n371), .Y(n472) );
  MUX2X1 U410 ( .B(n814), .A(n823), .S(n370), .Y(n488) );
  MUX2X1 U411 ( .B(n756), .A(n753), .S(n434), .Y(n1195) );
  MUX2X1 U412 ( .B(n756), .A(n757), .S(n368), .Y(n1163) );
  MUX2X1 U413 ( .B(n736), .A(n732), .S(n434), .Y(n1194) );
  MUX2X1 U414 ( .B(n736), .A(n1333), .S(n437), .Y(n1178) );
  MUX2X1 U415 ( .B(n736), .A(n735), .S(n368), .Y(n1162) );
  MUX2X1 U416 ( .B(n736), .A(n748), .S(n435), .Y(n1146) );
  MUX2X1 U417 ( .B(n736), .A(n734), .S(n369), .Y(n459) );
  MUX2X1 U418 ( .B(n329), .A(n733), .S(n370), .Y(n491) );
  MUX2X1 U419 ( .B(n329), .A(n1334), .S(n371), .Y(n475) );
  MUX2X1 U420 ( .B(n904), .A(n912), .S(n434), .Y(n1201) );
  MUX2X1 U421 ( .B(n904), .A(n913), .S(n437), .Y(n1185) );
  MUX2X1 U422 ( .B(n904), .A(n900), .S(n368), .Y(n1169) );
  INVX2 U423 ( .A(n525), .Y(n368) );
  MUX2X1 U424 ( .B(n904), .A(n901), .S(n435), .Y(n1153) );
  MUX2X1 U425 ( .B(n904), .A(n903), .S(n369), .Y(n452) );
  MUX2X1 U426 ( .B(n904), .A(n902), .S(n371), .Y(n468) );
  MUX2X1 U427 ( .B(n904), .A(n911), .S(n370), .Y(n484) );
  MUX2X1 U428 ( .B(n904), .A(n910), .S(n372), .Y(n500) );
  INVX8 U429 ( .A(w_data[4]), .Y(n715) );
  MUX2X1 U430 ( .B(n838), .A(n833), .S(n434), .Y(n1198) );
  MUX2X1 U431 ( .B(n838), .A(n1421), .S(n437), .Y(n1182) );
  MUX2X1 U432 ( .B(n838), .A(n848), .S(n435), .Y(n1150) );
  MUX2X1 U433 ( .B(n838), .A(n847), .S(n369), .Y(n455) );
  MUX2X1 U434 ( .B(n838), .A(n846), .S(n371), .Y(n471) );
  MUX2X1 U435 ( .B(n838), .A(n834), .S(n370), .Y(n487) );
  MUX2X1 U436 ( .B(n331), .A(n1418), .S(n372), .Y(n503) );
  MUX2X1 U437 ( .B(n331), .A(n1419), .S(n368), .Y(n1166) );
  INVX8 U438 ( .A(w_data[3]), .Y(n693) );
  MUX2X1 U439 ( .B(n883), .A(n1464), .S(n372), .Y(n501) );
  MUX2X1 U440 ( .B(n861), .A(n855), .S(n434), .Y(n1199) );
  MUX2X1 U441 ( .B(n861), .A(n856), .S(n437), .Y(n1183) );
  MUX2X1 U442 ( .B(n861), .A(n1444), .S(n368), .Y(n1167) );
  MUX2X1 U443 ( .B(n861), .A(n872), .S(n435), .Y(n1151) );
  MUX2X1 U444 ( .B(n861), .A(n870), .S(n369), .Y(n454) );
  MUX2X1 U445 ( .B(n861), .A(n857), .S(n370), .Y(n486) );
  MUX2X1 U446 ( .B(n861), .A(n1442), .S(n600), .Y(n502) );
  MUX2X1 U447 ( .B(n861), .A(n1441), .S(n371), .Y(n470) );
  INVX8 U448 ( .A(w_data[2]), .Y(n674) );
  MUX2X1 U449 ( .B(n946), .A(n954), .S(n434), .Y(n1203) );
  MUX2X1 U450 ( .B(n946), .A(n955), .S(n437), .Y(n1187) );
  MUX2X1 U451 ( .B(n946), .A(n942), .S(n368), .Y(n1171) );
  MUX2X1 U452 ( .B(n946), .A(n943), .S(n435), .Y(n1155) );
  MUX2X1 U453 ( .B(n946), .A(n945), .S(n609), .Y(n450) );
  MUX2X1 U454 ( .B(n946), .A(n944), .S(n607), .Y(n466) );
  MUX2X1 U455 ( .B(n946), .A(n953), .S(n605), .Y(n482) );
  MUX2X1 U456 ( .B(n946), .A(n952), .S(n372), .Y(n498) );
  MUX2X1 U457 ( .B(n925), .A(n921), .S(n368), .Y(n1170) );
  NAND2X1 U458 ( .A(n426), .B(n515), .Y(n373) );
  MUX2X1 U459 ( .B(n883), .A(n1476), .S(n434), .Y(n1200) );
  MUX2X1 U460 ( .B(n883), .A(n1467), .S(n437), .Y(n1184) );
  MUX2X1 U461 ( .B(n883), .A(n1474), .S(n368), .Y(n1168) );
  MUX2X1 U462 ( .B(n326), .A(n1466), .S(n435), .Y(n1152) );
  MUX2X1 U463 ( .B(n326), .A(n1472), .S(n609), .Y(n453) );
  MUX2X1 U464 ( .B(n332), .A(n1465), .S(n607), .Y(n469) );
  INVX1 U465 ( .A(r2_sel[1]), .Y(n374) );
  BUFX4 U466 ( .A(r2_sel[1]), .Y(n375) );
  BUFX4 U467 ( .A(n821), .Y(n376) );
  BUFX2 U468 ( .A(n1443), .Y(n377) );
  INVX1 U469 ( .A(n358), .Y(n845) );
  OAI22X1 U470 ( .A(n373), .B(n872), .C(n1444), .D(n871), .Y(n873) );
  NAND2X1 U471 ( .A(n379), .B(n378), .Y(r2_data[1]) );
  INVX1 U472 ( .A(n667), .Y(n378) );
  INVX1 U473 ( .A(n666), .Y(n379) );
  AND2X2 U474 ( .A(n821), .B(r2_sel[0]), .Y(n442) );
  NAND3X1 U475 ( .A(n362), .B(n381), .C(n380), .Y(r2_data[5]) );
  INVX1 U476 ( .A(n750), .Y(n380) );
  INVX2 U477 ( .A(n749), .Y(n381) );
  INVX1 U478 ( .A(n996), .Y(n552) );
  INVX4 U479 ( .A(r1_sel[1]), .Y(n1438) );
  INVX1 U480 ( .A(r2_sel[0]), .Y(n382) );
  INVX4 U481 ( .A(r2_sel[0]), .Y(n820) );
  INVX1 U482 ( .A(n397), .Y(n383) );
  INVX2 U483 ( .A(n801), .Y(n397) );
  INVX1 U484 ( .A(n1132), .Y(n384) );
  INVX1 U485 ( .A(n1074), .Y(n385) );
  NAND2X1 U486 ( .A(n851), .B(n386), .Y(r2_data[9]) );
  NOR2X1 U487 ( .A(n387), .B(n854), .Y(n386) );
  NAND2X1 U488 ( .A(n853), .B(n852), .Y(n387) );
  BUFX2 U489 ( .A(n1543), .Y(n388) );
  INVX4 U490 ( .A(n392), .Y(n406) );
  INVX1 U491 ( .A(n396), .Y(n389) );
  BUFX2 U492 ( .A(r1_sel[1]), .Y(n390) );
  INVX1 U493 ( .A(n342), .Y(n416) );
  AND2X2 U494 ( .A(n438), .B(n426), .Y(n684) );
  NAND3X1 U495 ( .A(n375), .B(n630), .C(n382), .Y(n392) );
  INVX2 U496 ( .A(n564), .Y(n393) );
  BUFX2 U497 ( .A(r2_sel[0]), .Y(n394) );
  AND2X2 U498 ( .A(n400), .B(n517), .Y(n396) );
  INVX1 U499 ( .A(n414), .Y(n398) );
  AND2X2 U500 ( .A(n563), .B(n1131), .Y(n1134) );
  AND2X1 U501 ( .A(n374), .B(n820), .Y(n515) );
  AND2X2 U502 ( .A(n647), .B(n395), .Y(n400) );
  INVX1 U503 ( .A(n1438), .Y(n399) );
  BUFX2 U504 ( .A(n892), .Y(n402) );
  INVX4 U505 ( .A(n550), .Y(n403) );
  INVX4 U506 ( .A(n550), .Y(n551) );
  INVX2 U507 ( .A(n552), .Y(n553) );
  MUX2X1 U508 ( .B(n332), .A(n1470), .S(n605), .Y(n485) );
  INVX2 U509 ( .A(n564), .Y(n1315) );
  BUFX2 U510 ( .A(n542), .Y(n404) );
  INVX2 U511 ( .A(n1072), .Y(n405) );
  INVX2 U512 ( .A(n1072), .Y(n1375) );
  MUX2X1 U513 ( .B(n789), .A(n798), .S(n609), .Y(n457) );
  INVX2 U514 ( .A(n1109), .Y(n407) );
  INVX1 U515 ( .A(n1109), .Y(n1361) );
  INVX2 U516 ( .A(n443), .Y(n408) );
  INVX2 U517 ( .A(n445), .Y(n409) );
  INVX1 U518 ( .A(n407), .Y(n411) );
  INVX1 U519 ( .A(n442), .Y(n656) );
  AND2X2 U520 ( .A(n442), .B(n426), .Y(n445) );
  INVX4 U521 ( .A(n446), .Y(n447) );
  INVX1 U522 ( .A(n1560), .Y(n412) );
  INVX1 U523 ( .A(n395), .Y(n413) );
  BUFX2 U524 ( .A(n868), .Y(n414) );
  BUFX4 U525 ( .A(n1445), .Y(n415) );
  AND2X2 U526 ( .A(n339), .B(n820), .Y(n418) );
  BUFX2 U527 ( .A(n1443), .Y(n419) );
  NAND2X1 U528 ( .A(n420), .B(\regs[6][4] ), .Y(n421) );
  NAND2X1 U529 ( .A(n421), .B(n1308), .Y(n1310) );
  INVX1 U530 ( .A(n1422), .Y(n420) );
  BUFX2 U531 ( .A(n775), .Y(n423) );
  INVX2 U532 ( .A(n775), .Y(n884) );
  INVX2 U533 ( .A(n322), .Y(n424) );
  MUX2X1 U534 ( .B(n925), .A(n933), .S(n434), .Y(n1202) );
  INVX2 U535 ( .A(n522), .Y(n434) );
  MUX2X1 U536 ( .B(n925), .A(n934), .S(n437), .Y(n1186) );
  INVX4 U537 ( .A(n892), .Y(n758) );
  OR2X2 U538 ( .A(r1_sel[2]), .B(r1_sel[3]), .Y(n1072) );
  AND2X2 U539 ( .A(n647), .B(r2_sel[2]), .Y(n426) );
  AND2X2 U540 ( .A(n521), .B(n532), .Y(n427) );
  INVX4 U541 ( .A(n427), .Y(n892) );
  MUX2X1 U542 ( .B(n925), .A(n931), .S(n600), .Y(n499) );
  MUX2X1 U543 ( .B(n925), .A(n922), .S(n435), .Y(n1154) );
  INVX2 U544 ( .A(n524), .Y(n435) );
  MUX2X1 U545 ( .B(n925), .A(n924), .S(n609), .Y(n451) );
  MUX2X1 U546 ( .B(n925), .A(n923), .S(n607), .Y(n467) );
  MUX2X1 U547 ( .B(n925), .A(n932), .S(n605), .Y(n483) );
  MUX2X1 U548 ( .B(n974), .A(n990), .S(n600), .Y(n497) );
  AND2X2 U549 ( .A(r2_sel[2]), .B(n647), .Y(n533) );
  INVX4 U550 ( .A(n373), .Y(n988) );
  NAND2X1 U551 ( .A(n1312), .B(n364), .Y(r1_data[4]) );
  AND2X2 U552 ( .A(n405), .B(r1_sel[1]), .Y(n433) );
  MUX2X1 U553 ( .B(n789), .A(n783), .S(n434), .Y(n1196) );
  MUX2X1 U554 ( .B(n789), .A(n784), .S(n437), .Y(n1180) );
  INVX2 U555 ( .A(n523), .Y(n437) );
  MUX2X1 U556 ( .B(n789), .A(n800), .S(n368), .Y(n1164) );
  MUX2X1 U557 ( .B(n789), .A(n802), .S(n435), .Y(n1148) );
  OR2X2 U558 ( .A(n660), .B(n659), .Y(n436) );
  NAND2X1 U559 ( .A(n436), .B(n658), .Y(n661) );
  MUX2X1 U560 ( .B(n756), .A(n754), .S(n609), .Y(n458) );
  MUX2X1 U561 ( .B(n756), .A(n755), .S(n607), .Y(n474) );
  MUX2X1 U562 ( .B(n756), .A(n777), .S(n605), .Y(n490) );
  MUX2X1 U563 ( .B(n328), .A(n776), .S(n600), .Y(n506) );
  MUX2X1 U564 ( .B(n328), .A(n1340), .S(n437), .Y(n1179) );
  BUFX2 U565 ( .A(n1439), .Y(n439) );
  OR2X1 U566 ( .A(n664), .B(n403), .Y(n440) );
  NAND2X1 U567 ( .A(n440), .B(n663), .Y(n667) );
  INVX8 U568 ( .A(w_data[8]), .Y(n814) );
  AND2X2 U569 ( .A(n533), .B(n519), .Y(n514) );
  NAND2X1 U570 ( .A(n1560), .B(\regs[6][9] ), .Y(n441) );
  NAND2X1 U571 ( .A(n1420), .B(n441), .Y(n1423) );
  NAND2X1 U572 ( .A(n363), .B(n1425), .Y(r1_data[9]) );
  INVX1 U573 ( .A(n382), .Y(n443) );
  INVX1 U574 ( .A(n799), .Y(n444) );
  MUX2X1 U575 ( .B(n789), .A(n797), .S(n607), .Y(n473) );
  MUX2X1 U576 ( .B(n789), .A(n785), .S(n605), .Y(n489) );
  MUX2X1 U577 ( .B(n789), .A(n602), .S(n600), .Y(n505) );
  OR2X2 U578 ( .A(n563), .B(n1119), .Y(n1445) );
  INVX4 U579 ( .A(n563), .Y(n565) );
  INVX4 U580 ( .A(n1475), .Y(n446) );
  AND2X2 U581 ( .A(n533), .B(n442), .Y(n448) );
  AND2X2 U582 ( .A(n533), .B(n418), .Y(n513) );
  AND2X2 U583 ( .A(r1_sel[1]), .B(n537), .Y(n518) );
  AND2X2 U584 ( .A(n375), .B(n820), .Y(n517) );
  AND2X2 U585 ( .A(n375), .B(r2_sel[0]), .Y(n519) );
  AND2X2 U586 ( .A(n375), .B(r2_sel[0]), .Y(n521) );
  AND2X1 U587 ( .A(n344), .B(r1_sel[3]), .Y(n535) );
  AND2X1 U588 ( .A(n413), .B(r2_sel[3]), .Y(n536) );
  INVX2 U589 ( .A(n1554), .Y(n1458) );
  INVX2 U590 ( .A(n763), .Y(n977) );
  AND2X2 U591 ( .A(n426), .B(n521), .Y(n516) );
  INVX2 U592 ( .A(n1568), .Y(n1459) );
  INVX2 U593 ( .A(n759), .Y(n975) );
  INVX2 U594 ( .A(n761), .Y(n976) );
  INVX2 U595 ( .A(n1570), .Y(n1453) );
  INVX2 U596 ( .A(n765), .Y(n978) );
  INVX2 U597 ( .A(n526), .Y(n569) );
  INVX2 U598 ( .A(n527), .Y(n568) );
  INVX2 U599 ( .A(n528), .Y(n567) );
  INVX2 U600 ( .A(n529), .Y(n566) );
  INVX2 U601 ( .A(n561), .Y(n562) );
  INVX2 U602 ( .A(n557), .Y(n558) );
  INVX2 U603 ( .A(n559), .Y(n560) );
  INVX2 U604 ( .A(n555), .Y(n556) );
  AND2X2 U605 ( .A(n521), .B(n426), .Y(n520) );
  AND2X2 U606 ( .A(n338), .B(n359), .Y(n522) );
  AND2X2 U607 ( .A(n359), .B(n337), .Y(n523) );
  AND2X2 U608 ( .A(n360), .B(n337), .Y(n524) );
  AND2X2 U609 ( .A(n360), .B(n338), .Y(n525) );
  INVX2 U610 ( .A(n619), .Y(n973) );
  INVX2 U611 ( .A(n616), .Y(n972) );
  INVX2 U613 ( .A(n614), .Y(n971) );
  INVX2 U614 ( .A(n611), .Y(n970) );
  INVX2 U615 ( .A(n1564), .Y(n561) );
  INVX2 U616 ( .A(n1566), .Y(n557) );
  INVX2 U617 ( .A(n1550), .Y(n555) );
  INVX2 U618 ( .A(n1548), .Y(n559) );
  AND2X2 U619 ( .A(n360), .B(n993), .Y(n526) );
  AND2X2 U620 ( .A(n360), .B(n995), .Y(n527) );
  AND2X2 U621 ( .A(n995), .B(n359), .Y(n529) );
  INVX2 U622 ( .A(n548), .Y(n549) );
  INVX2 U623 ( .A(n981), .Y(n548) );
  INVX2 U624 ( .A(n545), .Y(n546) );
  INVX2 U625 ( .A(n979), .Y(n545) );
  INVX2 U626 ( .A(n543), .Y(n544) );
  INVX2 U627 ( .A(n980), .Y(n543) );
  INVX2 U628 ( .A(n366), .Y(n547) );
  AND2X2 U629 ( .A(n985), .B(n399), .Y(n530) );
  AND2X2 U630 ( .A(n769), .B(n438), .Y(n531) );
  AND2X2 U631 ( .A(n647), .B(n345), .Y(n532) );
  AND2X2 U632 ( .A(n647), .B(n351), .Y(n534) );
  BUFX2 U633 ( .A(n570), .Y(n578) );
  BUFX2 U634 ( .A(n570), .Y(n579) );
  BUFX2 U635 ( .A(n570), .Y(n580) );
  BUFX2 U636 ( .A(n571), .Y(n581) );
  BUFX2 U637 ( .A(n571), .Y(n582) );
  BUFX2 U638 ( .A(n571), .Y(n583) );
  BUFX2 U639 ( .A(n572), .Y(n584) );
  BUFX2 U640 ( .A(n572), .Y(n585) );
  BUFX2 U641 ( .A(n572), .Y(n586) );
  BUFX2 U642 ( .A(n573), .Y(n587) );
  BUFX2 U643 ( .A(n573), .Y(n588) );
  BUFX2 U644 ( .A(n573), .Y(n589) );
  BUFX2 U645 ( .A(n574), .Y(n590) );
  BUFX2 U646 ( .A(n574), .Y(n591) );
  BUFX2 U647 ( .A(n574), .Y(n592) );
  BUFX2 U648 ( .A(n575), .Y(n593) );
  BUFX2 U649 ( .A(n575), .Y(n594) );
  BUFX2 U650 ( .A(n575), .Y(n595) );
  BUFX2 U651 ( .A(n576), .Y(n596) );
  BUFX2 U652 ( .A(n576), .Y(n597) );
  BUFX2 U653 ( .A(n576), .Y(n598) );
  BUFX2 U654 ( .A(n577), .Y(n599) );
  BUFX2 U655 ( .A(n_reset), .Y(n577) );
  BUFX2 U656 ( .A(n_reset), .Y(n570) );
  BUFX2 U657 ( .A(n_reset), .Y(n571) );
  BUFX2 U658 ( .A(n_reset), .Y(n572) );
  BUFX2 U659 ( .A(n_reset), .Y(n573) );
  BUFX2 U660 ( .A(n_reset), .Y(n574) );
  BUFX2 U661 ( .A(n_reset), .Y(n575) );
  BUFX2 U662 ( .A(n_reset), .Y(n576) );
  INVX8 U663 ( .A(w_data[6]), .Y(n756) );
  AND2X2 U664 ( .A(n1071), .B(r1_sel[2]), .Y(n537) );
  NAND2X1 U665 ( .A(n533), .B(n519), .Y(n538) );
  NAND2X1 U666 ( .A(n325), .B(n519), .Y(n539) );
  AND2X2 U667 ( .A(n405), .B(r1_sel[1]), .Y(n540) );
  INVX4 U668 ( .A(n540), .Y(n1473) );
  AND2X2 U669 ( .A(n407), .B(n391), .Y(n541) );
  OR2X2 U670 ( .A(n1439), .B(r1_sel[1]), .Y(n1475) );
  OR2X1 U671 ( .A(n878), .B(n879), .Y(r2_data[10]) );
  OR2X1 U672 ( .A(n808), .B(n809), .Y(r2_data[7]) );
  INVX8 U673 ( .A(n403), .Y(n893) );
  INVX8 U674 ( .A(w_data[5]), .Y(n736) );
  AND2X2 U675 ( .A(n537), .B(r1_sel[1]), .Y(n542) );
  INVX4 U676 ( .A(n542), .Y(n1477) );
  INVX8 U677 ( .A(w_data[12]), .Y(n904) );
  INVX4 U678 ( .A(n1088), .Y(n1562) );
  INVX4 U679 ( .A(n1087), .Y(n1561) );
  INVX4 U680 ( .A(n1445), .Y(n1544) );
  INVX8 U681 ( .A(w_data[7]), .Y(n789) );
  INVX8 U682 ( .A(w_data[9]), .Y(n838) );
  INVX8 U683 ( .A(w_data[14]), .Y(n946) );
  INVX8 U684 ( .A(w_data[11]), .Y(n883) );
  INVX8 U685 ( .A(w_data[10]), .Y(n861) );
  INVX8 U686 ( .A(w_data[15]), .Y(n974) );
  INVX8 U687 ( .A(w_data[13]), .Y(n925) );
  INVX4 U688 ( .A(w_data[0]), .Y(n620) );
  INVX4 U689 ( .A(n1070), .Y(n1543) );
  INVX4 U690 ( .A(n1073), .Y(n1546) );
  INVX4 U691 ( .A(n1074), .Y(n1545) );
  INVX8 U692 ( .A(r1_sel[0]), .Y(n563) );
  INVX8 U693 ( .A(n563), .Y(n564) );
  INVX2 U694 ( .A(outreg_data[0]), .Y(n1085) );
  INVX2 U695 ( .A(w_sel[2]), .Y(n618) );
  INVX2 U696 ( .A(w_sel[0]), .Y(n1578) );
  INVX2 U697 ( .A(w_sel[1]), .Y(n613) );
  NAND3X1 U698 ( .A(n365), .B(n1578), .C(n613), .Y(n600) );
  MUX2X1 U699 ( .B(n1085), .A(n620), .S(n603), .Y(n512) );
  INVX2 U700 ( .A(outreg_data[1]), .Y(n1097) );
  MUX2X1 U701 ( .B(n1097), .A(n645), .S(n603), .Y(n511) );
  INVX2 U702 ( .A(outreg_data[2]), .Y(n687) );
  MUX2X1 U703 ( .B(n687), .A(n674), .S(n603), .Y(n510) );
  INVX2 U704 ( .A(outreg_data[3]), .Y(n1287) );
  MUX2X1 U705 ( .B(n1287), .A(n693), .S(n603), .Y(n509) );
  INVX2 U706 ( .A(outreg_data[4]), .Y(n1306) );
  MUX2X1 U707 ( .B(n1306), .A(n715), .S(n603), .Y(n508) );
  INVX2 U708 ( .A(outreg_data[5]), .Y(n601) );
  MUX2X1 U709 ( .B(n601), .A(n736), .S(n603), .Y(n507) );
  INVX2 U710 ( .A(outreg_data[6]), .Y(n776) );
  INVX2 U711 ( .A(outreg_data[7]), .Y(n602) );
  INVX2 U712 ( .A(outreg_data[8]), .Y(n822) );
  MUX2X1 U713 ( .B(n822), .A(n814), .S(n603), .Y(n504) );
  INVX2 U714 ( .A(outreg_data[9]), .Y(n1418) );
  INVX2 U715 ( .A(outreg_data[10]), .Y(n1442) );
  INVX2 U716 ( .A(outreg_data[11]), .Y(n1464) );
  INVX2 U717 ( .A(outreg_data[12]), .Y(n910) );
  INVX2 U718 ( .A(outreg_data[13]), .Y(n931) );
  INVX2 U719 ( .A(outreg_data[14]), .Y(n952) );
  INVX2 U720 ( .A(outreg_data[15]), .Y(n990) );
  INVX2 U721 ( .A(\regs[7][0] ), .Y(n604) );
  MUX2X1 U722 ( .B(n604), .A(n620), .S(n522), .Y(n1189) );
  INVX2 U723 ( .A(\regs[6][0] ), .Y(n1090) );
  MUX2X1 U724 ( .B(n1090), .A(n620), .S(n523), .Y(n1173) );
  INVX2 U725 ( .A(\regs[1][0] ), .Y(n629) );
  NAND3X1 U726 ( .A(n365), .B(w_sel[0]), .C(n613), .Y(n605) );
  MUX2X1 U727 ( .B(n629), .A(n620), .S(n969), .Y(n496) );
  INVX2 U728 ( .A(\regs[5][0] ), .Y(n1086) );
  MUX2X1 U729 ( .B(n1086), .A(n620), .S(n525), .Y(n1157) );
  INVX2 U730 ( .A(\regs[4][0] ), .Y(n606) );
  MUX2X1 U731 ( .B(n606), .A(n620), .S(n524), .Y(n1141) );
  INVX2 U732 ( .A(\regs[2][0] ), .Y(n608) );
  NAND3X1 U733 ( .A(w_sel[1]), .B(n1578), .C(n365), .Y(n607) );
  MUX2X1 U734 ( .B(n608), .A(n620), .S(n965), .Y(n480) );
  INVX2 U735 ( .A(\regs[3][0] ), .Y(n610) );
  NAND3X1 U736 ( .A(w_sel[1]), .B(w_sel[0]), .C(n365), .Y(n609) );
  MUX2X1 U737 ( .B(n610), .A(n620), .S(n967), .Y(n464) );
  INVX2 U738 ( .A(\regs[9][0] ), .Y(n612) );
  NAND3X1 U739 ( .A(n995), .B(n618), .C(n613), .Y(n611) );
  MUX2X1 U740 ( .B(n612), .A(n620), .S(n970), .Y(n1221) );
  INVX2 U741 ( .A(\regs[8][0] ), .Y(n615) );
  NAND3X1 U742 ( .A(n993), .B(n618), .C(n613), .Y(n614) );
  MUX2X1 U743 ( .B(n615), .A(n620), .S(n971), .Y(n1205) );
  INVX2 U744 ( .A(\regs[11][0] ), .Y(n617) );
  NAND3X1 U745 ( .A(n995), .B(w_sel[1]), .C(n618), .Y(n616) );
  MUX2X1 U746 ( .B(n617), .A(n620), .S(n972), .Y(n1253) );
  INVX2 U747 ( .A(\regs[10][0] ), .Y(n621) );
  NAND3X1 U748 ( .A(n993), .B(w_sel[1]), .C(n618), .Y(n619) );
  MUX2X1 U749 ( .B(n621), .A(n620), .S(n973), .Y(n1237) );
  INVX2 U750 ( .A(r2_sel[3]), .Y(n647) );
  AOI22X1 U751 ( .A(n988), .B(\regs[4][0] ), .C(n416), .D(\regs[2][0] ), .Y(
        n636) );
  NAND3X1 U752 ( .A(n769), .B(n443), .C(n376), .Y(n761) );
  NAND3X1 U753 ( .A(n769), .B(n376), .C(n408), .Y(n759) );
  AOI22X1 U754 ( .A(n976), .B(\regs[9][0] ), .C(n975), .D(\regs[8][0] ), .Y(
        n626) );
  NAND2X1 U755 ( .A(n531), .B(n443), .Y(n765) );
  NAND2X1 U756 ( .A(n531), .B(n408), .Y(n763) );
  AOI22X1 U757 ( .A(n978), .B(\regs[11][0] ), .C(n977), .D(\regs[10][0] ), .Y(
        n625) );
  INVX2 U758 ( .A(\regs[13][0] ), .Y(n1076) );
  NAND3X1 U759 ( .A(n536), .B(n443), .C(n376), .Y(n980) );
  INVX2 U760 ( .A(\regs[12][0] ), .Y(n1075) );
  NAND3X1 U761 ( .A(n536), .B(n376), .C(n408), .Y(n979) );
  OAI22X1 U762 ( .A(n1076), .B(n544), .C(n1075), .D(n546), .Y(n623) );
  INVX2 U763 ( .A(\regs[15][0] ), .Y(n1078) );
  INVX2 U764 ( .A(\regs[14][0] ), .Y(n1077) );
  NAND3X1 U765 ( .A(n536), .B(n438), .C(n408), .Y(n981) );
  OAI22X1 U766 ( .A(n1078), .B(n547), .C(n1077), .D(n549), .Y(n622) );
  NOR2X1 U767 ( .A(n623), .B(n622), .Y(n624) );
  NAND3X1 U768 ( .A(n626), .B(n625), .C(n624), .Y(n627) );
  AOI21X1 U769 ( .A(n758), .B(\regs[3][0] ), .C(n627), .Y(n635) );
  NAND2X1 U770 ( .A(n533), .B(n442), .Y(n871) );
  NOR2X1 U771 ( .A(r2_sel[3]), .B(r2_sel[2]), .Y(n628) );
  NAND3X1 U772 ( .A(n374), .B(r2_sel[0]), .C(n628), .Y(n991) );
  OAI22X1 U773 ( .A(n1086), .B(n871), .C(n629), .D(n430), .Y(n633) );
  NOR2X1 U774 ( .A(r2_sel[3]), .B(n351), .Y(n630) );
  NAND3X1 U775 ( .A(n375), .B(n820), .C(n630), .Y(n996) );
  NAND3X1 U776 ( .A(n376), .B(n820), .C(n534), .Y(n775) );
  AOI22X1 U777 ( .A(n520), .B(\regs[7][0] ), .C(outreg_data[0]), .D(n341), .Y(
        n631) );
  OAI21X1 U778 ( .A(n1090), .B(n553), .C(n631), .Y(n632) );
  NOR2X1 U779 ( .A(n633), .B(n632), .Y(n634) );
  NAND3X1 U780 ( .A(n636), .B(n635), .C(n634), .Y(r2_data[0]) );
  INVX2 U781 ( .A(\regs[7][1] ), .Y(n637) );
  MUX2X1 U782 ( .B(n637), .A(n645), .S(n522), .Y(n1190) );
  INVX2 U783 ( .A(\regs[6][1] ), .Y(n638) );
  MUX2X1 U784 ( .B(n638), .A(n645), .S(n523), .Y(n1174) );
  INVX2 U785 ( .A(\regs[1][1] ), .Y(n664) );
  MUX2X1 U786 ( .B(n664), .A(n645), .S(n969), .Y(n495) );
  INVX2 U787 ( .A(\regs[3][1] ), .Y(n639) );
  MUX2X1 U788 ( .B(n639), .A(n645), .S(n967), .Y(n463) );
  INVX2 U789 ( .A(\regs[2][1] ), .Y(n1096) );
  MUX2X1 U790 ( .B(n1096), .A(n645), .S(n965), .Y(n479) );
  INVX2 U791 ( .A(\regs[4][1] ), .Y(n640) );
  MUX2X1 U792 ( .B(n640), .A(n645), .S(n524), .Y(n1142) );
  INVX2 U793 ( .A(\regs[5][1] ), .Y(n641) );
  MUX2X1 U794 ( .B(n641), .A(n645), .S(n525), .Y(n1158) );
  INVX2 U795 ( .A(\regs[9][1] ), .Y(n642) );
  MUX2X1 U796 ( .B(n642), .A(n645), .S(n970), .Y(n1222) );
  INVX2 U797 ( .A(\regs[8][1] ), .Y(n643) );
  MUX2X1 U798 ( .B(n643), .A(n645), .S(n971), .Y(n1206) );
  INVX2 U799 ( .A(\regs[11][1] ), .Y(n644) );
  MUX2X1 U800 ( .B(n644), .A(n645), .S(n972), .Y(n1254) );
  INVX2 U801 ( .A(\regs[10][1] ), .Y(n646) );
  MUX2X1 U802 ( .B(n646), .A(n645), .S(n973), .Y(n1238) );
  NAND2X1 U803 ( .A(n533), .B(\regs[5][1] ), .Y(n655) );
  AOI22X1 U804 ( .A(n548), .B(\regs[14][1] ), .C(n366), .D(\regs[15][1] ), .Y(
        n649) );
  AOI22X1 U805 ( .A(n545), .B(\regs[12][1] ), .C(n543), .D(\regs[13][1] ), .Y(
        n648) );
  NAND2X1 U806 ( .A(n649), .B(n648), .Y(n653) );
  AOI22X1 U807 ( .A(n976), .B(\regs[9][1] ), .C(n975), .D(\regs[8][1] ), .Y(
        n651) );
  AOI22X1 U808 ( .A(n978), .B(\regs[11][1] ), .C(n977), .D(\regs[10][1] ), .Y(
        n650) );
  NAND2X1 U809 ( .A(n651), .B(n650), .Y(n652) );
  NOR2X1 U810 ( .A(n653), .B(n652), .Y(n654) );
  OAI21X1 U811 ( .A(n656), .B(n655), .C(n654), .Y(n662) );
  OAI21X1 U812 ( .A(\regs[2][1] ), .B(n394), .C(n438), .Y(n660) );
  NOR2X1 U814 ( .A(n346), .B(r2_sel[3]), .Y(n657) );
  OAI21X1 U815 ( .A(\regs[3][1] ), .B(n382), .C(n657), .Y(n659) );
  NAND3X1 U816 ( .A(n418), .B(n325), .C(\regs[4][1] ), .Y(n658) );
  NOR2X1 U817 ( .A(n662), .B(n661), .Y(n663) );
  AOI22X1 U818 ( .A(n520), .B(\regs[7][1] ), .C(n406), .D(\regs[6][1] ), .Y(
        n665) );
  OAI21X1 U819 ( .A(n1097), .B(n423), .C(n665), .Y(n666) );
  INVX2 U820 ( .A(\regs[7][2] ), .Y(n1120) );
  MUX2X1 U821 ( .B(n1120), .A(n674), .S(n522), .Y(n1191) );
  INVX2 U822 ( .A(\regs[6][2] ), .Y(n683) );
  MUX2X1 U823 ( .B(n683), .A(n674), .S(n523), .Y(n1175) );
  INVX2 U824 ( .A(\regs[1][2] ), .Y(n682) );
  MUX2X1 U825 ( .B(n682), .A(n674), .S(n969), .Y(n494) );
  INVX2 U826 ( .A(\regs[5][2] ), .Y(n1118) );
  MUX2X1 U827 ( .B(n1118), .A(n674), .S(n525), .Y(n1159) );
  INVX2 U828 ( .A(\regs[4][2] ), .Y(n668) );
  MUX2X1 U829 ( .B(n668), .A(n674), .S(n524), .Y(n1143) );
  INVX2 U830 ( .A(\regs[2][2] ), .Y(n669) );
  MUX2X1 U831 ( .B(n669), .A(n674), .S(n965), .Y(n478) );
  INVX2 U832 ( .A(\regs[3][2] ), .Y(n670) );
  MUX2X1 U833 ( .B(n670), .A(n674), .S(n967), .Y(n462) );
  INVX2 U834 ( .A(\regs[9][2] ), .Y(n671) );
  MUX2X1 U835 ( .B(n671), .A(n674), .S(n970), .Y(n1223) );
  INVX2 U836 ( .A(\regs[8][2] ), .Y(n672) );
  MUX2X1 U837 ( .B(n672), .A(n674), .S(n971), .Y(n1207) );
  INVX2 U838 ( .A(\regs[11][2] ), .Y(n673) );
  MUX2X1 U839 ( .B(n673), .A(n674), .S(n972), .Y(n1255) );
  INVX2 U840 ( .A(\regs[10][2] ), .Y(n675) );
  MUX2X1 U841 ( .B(n675), .A(n674), .S(n973), .Y(n1239) );
  NAND2X1 U842 ( .A(n533), .B(n418), .Y(n801) );
  AOI22X1 U843 ( .A(n513), .B(\regs[4][2] ), .C(n432), .D(\regs[2][2] ), .Y(
        n692) );
  AOI22X1 U844 ( .A(n976), .B(\regs[9][2] ), .C(n975), .D(\regs[8][2] ), .Y(
        n680) );
  AOI22X1 U845 ( .A(n978), .B(\regs[11][2] ), .C(n977), .D(\regs[10][2] ), .Y(
        n679) );
  INVX2 U846 ( .A(\regs[13][2] ), .Y(n1122) );
  INVX2 U847 ( .A(\regs[12][2] ), .Y(n1121) );
  OAI22X1 U848 ( .A(n1122), .B(n544), .C(n1121), .D(n546), .Y(n677) );
  INVX2 U849 ( .A(\regs[15][2] ), .Y(n1124) );
  INVX2 U850 ( .A(\regs[14][2] ), .Y(n1123) );
  OAI22X1 U851 ( .A(n1124), .B(n547), .C(n1123), .D(n549), .Y(n676) );
  NOR2X1 U852 ( .A(n677), .B(n676), .Y(n678) );
  NAND3X1 U853 ( .A(n680), .B(n679), .C(n678), .Y(n681) );
  AOI21X1 U854 ( .A(n349), .B(\regs[3][2] ), .C(n681), .Y(n691) );
  NAND2X1 U855 ( .A(n426), .B(n442), .Y(n799) );
  OAI22X1 U856 ( .A(n1118), .B(n799), .C(n682), .D(n551), .Y(n689) );
  NOR2X1 U857 ( .A(n394), .B(n683), .Y(n685) );
  AOI22X1 U858 ( .A(n516), .B(\regs[7][2] ), .C(n685), .D(n684), .Y(n686) );
  OAI21X1 U859 ( .A(n775), .B(n687), .C(n686), .Y(n688) );
  NOR2X1 U860 ( .A(n689), .B(n688), .Y(n690) );
  NAND3X1 U861 ( .A(n692), .B(n691), .C(n690), .Y(r2_data[2]) );
  INVX2 U862 ( .A(\regs[4][3] ), .Y(n1285) );
  MUX2X1 U863 ( .B(n1285), .A(n693), .S(n524), .Y(n1144) );
  INVX2 U864 ( .A(\regs[2][3] ), .Y(n1288) );
  MUX2X1 U865 ( .B(n1288), .A(n693), .S(n965), .Y(n477) );
  INVX2 U866 ( .A(\regs[3][3] ), .Y(n1273) );
  MUX2X1 U867 ( .B(n1273), .A(n693), .S(n967), .Y(n461) );
  INVX2 U868 ( .A(\regs[6][3] ), .Y(n1286) );
  MUX2X1 U869 ( .B(n1286), .A(n693), .S(n523), .Y(n1176) );
  INVX2 U870 ( .A(\regs[1][3] ), .Y(n1272) );
  MUX2X1 U871 ( .B(n1272), .A(n693), .S(n969), .Y(n493) );
  INVX2 U872 ( .A(\regs[7][3] ), .Y(n1271) );
  MUX2X1 U873 ( .B(n1271), .A(n693), .S(n522), .Y(n1192) );
  INVX2 U874 ( .A(\regs[5][3] ), .Y(n1270) );
  MUX2X1 U875 ( .B(n1270), .A(n693), .S(n525), .Y(n1160) );
  INVX2 U876 ( .A(\regs[10][3] ), .Y(n698) );
  MUX2X1 U877 ( .B(n698), .A(n693), .S(n973), .Y(n1240) );
  INVX2 U878 ( .A(\regs[11][3] ), .Y(n699) );
  MUX2X1 U879 ( .B(n699), .A(n693), .S(n972), .Y(n1256) );
  INVX2 U880 ( .A(\regs[8][3] ), .Y(n696) );
  MUX2X1 U881 ( .B(n696), .A(n693), .S(n971), .Y(n1208) );
  INVX2 U882 ( .A(\regs[9][3] ), .Y(n697) );
  MUX2X1 U883 ( .B(n697), .A(n693), .S(n970), .Y(n1224) );
  AOI22X1 U884 ( .A(n355), .B(\regs[4][3] ), .C(n422), .D(outreg_data[3]), .Y(
        n709) );
  AOI22X1 U885 ( .A(n401), .B(\regs[2][3] ), .C(n758), .D(\regs[3][3] ), .Y(
        n708) );
  INVX2 U886 ( .A(\regs[14][3] ), .Y(n1278) );
  INVX2 U887 ( .A(\regs[15][3] ), .Y(n1279) );
  OAI22X1 U888 ( .A(n1278), .B(n549), .C(n1279), .D(n547), .Y(n695) );
  INVX2 U889 ( .A(\regs[12][3] ), .Y(n1276) );
  INVX2 U890 ( .A(\regs[13][3] ), .Y(n1277) );
  OAI22X1 U891 ( .A(n1276), .B(n546), .C(n1277), .D(n544), .Y(n694) );
  NOR2X1 U892 ( .A(n695), .B(n694), .Y(n704) );
  OAI22X1 U893 ( .A(n697), .B(n761), .C(n696), .D(n759), .Y(n701) );
  OAI22X1 U894 ( .A(n699), .B(n765), .C(n698), .D(n763), .Y(n700) );
  NOR2X1 U895 ( .A(n701), .B(n700), .Y(n703) );
  AOI22X1 U896 ( .A(n520), .B(\regs[7][3] ), .C(n445), .D(\regs[5][3] ), .Y(
        n702) );
  NAND3X1 U897 ( .A(n704), .B(n703), .C(n702), .Y(n706) );
  OAI22X1 U898 ( .A(n1272), .B(n551), .C(n322), .D(n1286), .Y(n705) );
  NOR2X1 U899 ( .A(n706), .B(n705), .Y(n707) );
  NAND3X1 U900 ( .A(n707), .B(n709), .C(n708), .Y(r2_data[3]) );
  INVX2 U901 ( .A(\regs[7][4] ), .Y(n710) );
  MUX2X1 U902 ( .B(n710), .A(n715), .S(n522), .Y(n1193) );
  INVX2 U903 ( .A(\regs[6][4] ), .Y(n1309) );
  MUX2X1 U904 ( .B(n1309), .A(n715), .S(n523), .Y(n1177) );
  INVX2 U905 ( .A(\regs[1][4] ), .Y(n711) );
  MUX2X1 U906 ( .B(n711), .A(n715), .S(n969), .Y(n492) );
  INVX2 U907 ( .A(\regs[5][4] ), .Y(n1307) );
  MUX2X1 U908 ( .B(n1307), .A(n715), .S(n525), .Y(n1161) );
  INVX2 U909 ( .A(\regs[4][4] ), .Y(n724) );
  MUX2X1 U910 ( .B(n724), .A(n715), .S(n524), .Y(n1145) );
  INVX2 U911 ( .A(\regs[2][4] ), .Y(n722) );
  MUX2X1 U912 ( .B(n722), .A(n715), .S(n965), .Y(n476) );
  INVX2 U913 ( .A(\regs[3][4] ), .Y(n723) );
  MUX2X1 U914 ( .B(n723), .A(n715), .S(n967), .Y(n460) );
  INVX2 U915 ( .A(\regs[9][4] ), .Y(n712) );
  MUX2X1 U916 ( .B(n712), .A(n367), .S(n970), .Y(n1225) );
  INVX2 U917 ( .A(\regs[8][4] ), .Y(n713) );
  MUX2X1 U918 ( .B(n713), .A(n715), .S(n971), .Y(n1209) );
  INVX2 U919 ( .A(\regs[11][4] ), .Y(n714) );
  MUX2X1 U920 ( .B(n714), .A(n367), .S(n972), .Y(n1257) );
  INVX2 U921 ( .A(\regs[10][4] ), .Y(n716) );
  MUX2X1 U922 ( .B(n716), .A(n715), .S(n973), .Y(n1241) );
  AOI22X1 U923 ( .A(n976), .B(\regs[9][4] ), .C(n975), .D(\regs[8][4] ), .Y(
        n721) );
  AOI22X1 U924 ( .A(n978), .B(\regs[11][4] ), .C(n977), .D(\regs[10][4] ), .Y(
        n720) );
  INVX2 U925 ( .A(\regs[13][4] ), .Y(n1297) );
  INVX2 U926 ( .A(\regs[12][4] ), .Y(n1296) );
  OAI22X1 U927 ( .A(n1297), .B(n544), .C(n1296), .D(n546), .Y(n718) );
  INVX2 U928 ( .A(\regs[15][4] ), .Y(n1299) );
  INVX2 U929 ( .A(\regs[14][4] ), .Y(n1298) );
  OAI22X1 U930 ( .A(n1299), .B(n547), .C(n1298), .D(n549), .Y(n717) );
  NOR2X1 U931 ( .A(n718), .B(n717), .Y(n719) );
  NAND3X1 U932 ( .A(n721), .B(n720), .C(n719), .Y(n731) );
  AOI22X1 U933 ( .A(n352), .B(\regs[7][4] ), .C(n348), .D(outreg_data[4]), .Y(
        n729) );
  AOI22X1 U934 ( .A(n424), .B(\regs[6][4] ), .C(n893), .D(\regs[1][4] ), .Y(
        n728) );
  OAI22X1 U935 ( .A(n723), .B(n402), .C(n722), .D(n389), .Y(n726) );
  OAI22X1 U936 ( .A(n724), .B(n425), .C(n1307), .D(n409), .Y(n725) );
  NOR2X1 U937 ( .A(n726), .B(n725), .Y(n727) );
  NAND3X1 U938 ( .A(n729), .B(n728), .C(n727), .Y(n730) );
  OR2X2 U939 ( .A(n731), .B(n730), .Y(r2_data[4]) );
  INVX2 U940 ( .A(\regs[7][5] ), .Y(n732) );
  INVX2 U941 ( .A(\regs[1][5] ), .Y(n733) );
  INVX2 U942 ( .A(\regs[6][5] ), .Y(n1333) );
  INVX2 U943 ( .A(\regs[3][5] ), .Y(n734) );
  INVX2 U944 ( .A(\regs[2][5] ), .Y(n1334) );
  INVX2 U945 ( .A(\regs[4][5] ), .Y(n748) );
  INVX2 U946 ( .A(\regs[5][5] ), .Y(n735) );
  INVX2 U947 ( .A(\regs[10][5] ), .Y(n741) );
  MUX2X1 U948 ( .B(n741), .A(n736), .S(n973), .Y(n1242) );
  INVX2 U949 ( .A(\regs[11][5] ), .Y(n742) );
  MUX2X1 U950 ( .B(n742), .A(n736), .S(n972), .Y(n1258) );
  INVX2 U951 ( .A(\regs[8][5] ), .Y(n739) );
  MUX2X1 U952 ( .B(n739), .A(n736), .S(n971), .Y(n1210) );
  INVX2 U953 ( .A(\regs[9][5] ), .Y(n740) );
  MUX2X1 U954 ( .B(n740), .A(n736), .S(n970), .Y(n1226) );
  AOI22X1 U955 ( .A(n514), .B(\regs[7][5] ), .C(n893), .D(\regs[1][5] ), .Y(
        n752) );
  AOI22X1 U956 ( .A(n406), .B(\regs[6][5] ), .C(\regs[3][5] ), .D(n758), .Y(
        n751) );
  INVX2 U957 ( .A(\regs[14][5] ), .Y(n1323) );
  INVX2 U958 ( .A(\regs[15][5] ), .Y(n1324) );
  OAI22X1 U959 ( .A(n1323), .B(n549), .C(n1324), .D(n547), .Y(n738) );
  INVX2 U960 ( .A(\regs[12][5] ), .Y(n1321) );
  INVX2 U961 ( .A(\regs[13][5] ), .Y(n1322) );
  OAI22X1 U962 ( .A(n1321), .B(n546), .C(n1322), .D(n544), .Y(n737) );
  NOR2X1 U963 ( .A(n738), .B(n737), .Y(n747) );
  OAI22X1 U964 ( .A(n740), .B(n761), .C(n739), .D(n759), .Y(n744) );
  OAI22X1 U965 ( .A(n742), .B(n765), .C(n741), .D(n763), .Y(n743) );
  NOR2X1 U966 ( .A(n744), .B(n743), .Y(n746) );
  AOI22X1 U967 ( .A(n445), .B(\regs[5][5] ), .C(outreg_data[5]), .D(n884), .Y(
        n745) );
  NAND3X1 U968 ( .A(n747), .B(n746), .C(n745), .Y(n750) );
  OAI22X1 U969 ( .A(n748), .B(n383), .C(n1334), .D(n389), .Y(n749) );
  INVX2 U970 ( .A(\regs[1][6] ), .Y(n777) );
  INVX2 U971 ( .A(\regs[10][6] ), .Y(n764) );
  MUX2X1 U972 ( .B(n764), .A(n756), .S(n973), .Y(n1243) );
  INVX2 U973 ( .A(\regs[11][6] ), .Y(n766) );
  MUX2X1 U974 ( .B(n766), .A(n756), .S(n972), .Y(n1259) );
  INVX2 U975 ( .A(\regs[8][6] ), .Y(n760) );
  MUX2X1 U976 ( .B(n760), .A(n756), .S(n971), .Y(n1211) );
  INVX2 U977 ( .A(\regs[9][6] ), .Y(n762) );
  MUX2X1 U978 ( .B(n762), .A(n756), .S(n970), .Y(n1227) );
  INVX2 U979 ( .A(\regs[7][6] ), .Y(n753) );
  INVX2 U980 ( .A(\regs[6][6] ), .Y(n1340) );
  INVX2 U981 ( .A(\regs[3][6] ), .Y(n754) );
  INVX2 U982 ( .A(\regs[2][6] ), .Y(n755) );
  INVX2 U983 ( .A(\regs[4][6] ), .Y(n1341) );
  MUX2X1 U984 ( .B(n1341), .A(n756), .S(n524), .Y(n1147) );
  INVX2 U985 ( .A(\regs[5][6] ), .Y(n757) );
  AOI22X1 U986 ( .A(\regs[3][6] ), .B(n758), .C(n356), .D(\regs[2][6] ), .Y(
        n782) );
  AOI22X1 U987 ( .A(n397), .B(\regs[4][6] ), .C(n444), .D(\regs[5][6] ), .Y(
        n781) );
  AOI22X1 U988 ( .A(n543), .B(\regs[13][6] ), .C(n545), .D(\regs[12][6] ), .Y(
        n772) );
  AOI22X1 U989 ( .A(n366), .B(\regs[15][6] ), .C(n548), .D(\regs[14][6] ), .Y(
        n771) );
  OAI22X1 U990 ( .A(n762), .B(n761), .C(n760), .D(n759), .Y(n768) );
  OAI22X1 U991 ( .A(n766), .B(n765), .C(n764), .D(n763), .Y(n767) );
  NOR2X1 U992 ( .A(n768), .B(n767), .Y(n770) );
  NAND3X1 U993 ( .A(n772), .B(n771), .C(n770), .Y(n773) );
  AOI21X1 U994 ( .A(n516), .B(\regs[7][6] ), .C(n773), .Y(n774) );
  OAI21X1 U995 ( .A(n1340), .B(n322), .C(n774), .Y(n779) );
  OAI22X1 U996 ( .A(n777), .B(n551), .C(n776), .D(n429), .Y(n778) );
  NOR2X1 U997 ( .A(n779), .B(n778), .Y(n780) );
  NAND3X1 U998 ( .A(n781), .B(n782), .C(n780), .Y(r2_data[6]) );
  INVX2 U999 ( .A(\regs[7][7] ), .Y(n783) );
  INVX2 U1000 ( .A(\regs[6][7] ), .Y(n784) );
  INVX2 U1001 ( .A(\regs[1][7] ), .Y(n785) );
  INVX2 U1002 ( .A(\regs[5][7] ), .Y(n800) );
  INVX2 U1003 ( .A(\regs[4][7] ), .Y(n802) );
  INVX2 U1004 ( .A(\regs[2][7] ), .Y(n797) );
  INVX2 U1005 ( .A(\regs[3][7] ), .Y(n798) );
  INVX2 U1006 ( .A(\regs[9][7] ), .Y(n786) );
  MUX2X1 U1007 ( .B(n786), .A(n431), .S(n970), .Y(n1228) );
  INVX2 U1008 ( .A(\regs[8][7] ), .Y(n787) );
  MUX2X1 U1009 ( .B(n787), .A(n431), .S(n971), .Y(n1212) );
  INVX2 U1010 ( .A(\regs[11][7] ), .Y(n788) );
  MUX2X1 U1011 ( .B(n788), .A(n431), .S(n972), .Y(n1260) );
  INVX2 U1012 ( .A(\regs[10][7] ), .Y(n790) );
  MUX2X1 U1013 ( .B(n790), .A(n431), .S(n973), .Y(n1244) );
  AOI22X1 U1014 ( .A(n976), .B(\regs[9][7] ), .C(n975), .D(\regs[8][7] ), .Y(
        n795) );
  AOI22X1 U1015 ( .A(n978), .B(\regs[11][7] ), .C(n977), .D(\regs[10][7] ), 
        .Y(n794) );
  INVX2 U1016 ( .A(\regs[13][7] ), .Y(n1367) );
  INVX2 U1017 ( .A(\regs[12][7] ), .Y(n1366) );
  OAI22X1 U1018 ( .A(n1367), .B(n544), .C(n1366), .D(n546), .Y(n792) );
  INVX2 U1020 ( .A(\regs[15][7] ), .Y(n1369) );
  INVX2 U1021 ( .A(\regs[14][7] ), .Y(n1368) );
  OAI22X1 U1022 ( .A(n1369), .B(n547), .C(n1368), .D(n549), .Y(n791) );
  NOR2X1 U1023 ( .A(n792), .B(n791), .Y(n793) );
  NAND3X1 U1024 ( .A(n795), .B(n794), .C(n793), .Y(n809) );
  AOI22X1 U1025 ( .A(n514), .B(\regs[7][7] ), .C(outreg_data[7]), .D(n884), 
        .Y(n807) );
  AOI22X1 U1026 ( .A(\regs[6][7] ), .B(n406), .C(n357), .D(\regs[1][7] ), .Y(
        n806) );
  OAI22X1 U1027 ( .A(n798), .B(n892), .C(n797), .D(n796), .Y(n804) );
  OAI22X1 U1028 ( .A(n802), .B(n801), .C(n800), .D(n799), .Y(n803) );
  NOR2X1 U1029 ( .A(n803), .B(n804), .Y(n805) );
  NAND3X1 U1030 ( .A(n807), .B(n806), .C(n805), .Y(n808) );
  INVX2 U1031 ( .A(\regs[5][8] ), .Y(n810) );
  INVX2 U1032 ( .A(\regs[4][8] ), .Y(n811) );
  INVX2 U1033 ( .A(\regs[2][8] ), .Y(n812) );
  INVX2 U1034 ( .A(\regs[3][8] ), .Y(n813) );
  INVX2 U1035 ( .A(\regs[7][8] ), .Y(n824) );
  INVX2 U1036 ( .A(\regs[6][8] ), .Y(n825) );
  INVX2 U1037 ( .A(\regs[1][8] ), .Y(n823) );
  INVX2 U1038 ( .A(\regs[9][8] ), .Y(n1390) );
  MUX2X1 U1039 ( .B(n1390), .A(n327), .S(n970), .Y(n1229) );
  INVX2 U1040 ( .A(\regs[8][8] ), .Y(n1399) );
  MUX2X1 U1041 ( .B(n1399), .A(n327), .S(n971), .Y(n1213) );
  INVX2 U1042 ( .A(\regs[11][8] ), .Y(n1391) );
  MUX2X1 U1043 ( .B(n1391), .A(n327), .S(n972), .Y(n1261) );
  INVX2 U1044 ( .A(\regs[10][8] ), .Y(n1400) );
  MUX2X1 U1045 ( .B(n1400), .A(n327), .S(n973), .Y(n1245) );
  AOI22X1 U1046 ( .A(n976), .B(\regs[9][8] ), .C(n975), .D(\regs[8][8] ), .Y(
        n819) );
  AOI22X1 U1047 ( .A(n978), .B(\regs[11][8] ), .C(n977), .D(\regs[10][8] ), 
        .Y(n818) );
  INVX2 U1048 ( .A(\regs[13][8] ), .Y(n1389) );
  INVX2 U1049 ( .A(\regs[12][8] ), .Y(n1398) );
  OAI22X1 U1050 ( .A(n1389), .B(n544), .C(n1398), .D(n546), .Y(n816) );
  INVX2 U1051 ( .A(\regs[15][8] ), .Y(n1388) );
  INVX2 U1052 ( .A(\regs[14][8] ), .Y(n1397) );
  OAI22X1 U1053 ( .A(n1388), .B(n547), .C(n1397), .D(n549), .Y(n815) );
  NOR2X1 U1054 ( .A(n816), .B(n815), .Y(n817) );
  NAND3X1 U1055 ( .A(n819), .B(n818), .C(n817), .Y(n832) );
  AOI22X1 U1056 ( .A(\regs[5][8] ), .B(n448), .C(\regs[4][8] ), .D(n988), .Y(
        n830) );
  NAND2X1 U1057 ( .A(n517), .B(n534), .Y(n868) );
  NAND2X1 U1058 ( .A(n519), .B(n400), .Y(n869) );
  AOI22X1 U1059 ( .A(n432), .B(\regs[2][8] ), .C(n410), .D(\regs[3][8] ), .Y(
        n829) );
  NAND3X1 U1060 ( .A(n376), .B(n820), .C(n532), .Y(n989) );
  OAI22X1 U1061 ( .A(n823), .B(n551), .C(n822), .D(n429), .Y(n827) );
  OAI22X1 U1062 ( .A(n322), .B(n825), .C(n824), .D(n538), .Y(n826) );
  NOR2X1 U1063 ( .A(n826), .B(n827), .Y(n828) );
  NAND3X1 U1064 ( .A(n830), .B(n829), .C(n828), .Y(n831) );
  INVX2 U1065 ( .A(\regs[7][9] ), .Y(n833) );
  INVX2 U1066 ( .A(\regs[6][9] ), .Y(n1421) );
  INVX2 U1067 ( .A(\regs[1][9] ), .Y(n834) );
  INVX2 U1068 ( .A(\regs[5][9] ), .Y(n1419) );
  INVX2 U1069 ( .A(\regs[4][9] ), .Y(n848) );
  INVX2 U1070 ( .A(\regs[2][9] ), .Y(n846) );
  INVX2 U1071 ( .A(\regs[3][9] ), .Y(n847) );
  INVX2 U1072 ( .A(\regs[9][9] ), .Y(n835) );
  MUX2X1 U1073 ( .B(n835), .A(n838), .S(n970), .Y(n1230) );
  INVX2 U1074 ( .A(\regs[8][9] ), .Y(n836) );
  MUX2X1 U1075 ( .B(n836), .A(n838), .S(n971), .Y(n1214) );
  INVX2 U1076 ( .A(\regs[11][9] ), .Y(n837) );
  MUX2X1 U1077 ( .B(n837), .A(n838), .S(n972), .Y(n1262) );
  INVX2 U1078 ( .A(\regs[10][9] ), .Y(n839) );
  MUX2X1 U1079 ( .B(n839), .A(n838), .S(n973), .Y(n1246) );
  AOI22X1 U1080 ( .A(n976), .B(\regs[9][9] ), .C(n975), .D(\regs[8][9] ), .Y(
        n844) );
  AOI22X1 U1081 ( .A(n978), .B(\regs[11][9] ), .C(n977), .D(\regs[10][9] ), 
        .Y(n843) );
  INVX2 U1082 ( .A(\regs[13][9] ), .Y(n1409) );
  INVX2 U1083 ( .A(\regs[12][9] ), .Y(n1408) );
  OAI22X1 U1084 ( .A(n1409), .B(n544), .C(n1408), .D(n546), .Y(n841) );
  INVX2 U1085 ( .A(\regs[15][9] ), .Y(n1411) );
  INVX2 U1086 ( .A(\regs[14][9] ), .Y(n1410) );
  OAI22X1 U1087 ( .A(n1411), .B(n547), .C(n1410), .D(n549), .Y(n840) );
  NOR2X1 U1088 ( .A(n841), .B(n840), .Y(n842) );
  NAND3X1 U1089 ( .A(n844), .B(n843), .C(n842), .Y(n854) );
  AOI22X1 U1090 ( .A(n514), .B(\regs[7][9] ), .C(n845), .D(outreg_data[9]), 
        .Y(n853) );
  AOI22X1 U1091 ( .A(n406), .B(\regs[6][9] ), .C(n357), .D(\regs[1][9] ), .Y(
        n852) );
  OAI22X1 U1092 ( .A(n847), .B(n340), .C(n846), .D(n414), .Y(n850) );
  OAI22X1 U1093 ( .A(n425), .B(n848), .C(n1419), .D(n409), .Y(n849) );
  NOR2X1 U1094 ( .A(n849), .B(n850), .Y(n851) );
  INVX2 U1095 ( .A(\regs[7][10] ), .Y(n855) );
  INVX2 U1096 ( .A(\regs[6][10] ), .Y(n856) );
  INVX2 U1097 ( .A(\regs[1][10] ), .Y(n857) );
  INVX2 U1098 ( .A(\regs[4][10] ), .Y(n872) );
  INVX2 U1099 ( .A(\regs[2][10] ), .Y(n1441) );
  INVX2 U1100 ( .A(\regs[3][10] ), .Y(n870) );
  INVX2 U1101 ( .A(\regs[9][10] ), .Y(n858) );
  MUX2X1 U1102 ( .B(n858), .A(n334), .S(n970), .Y(n1231) );
  INVX2 U1103 ( .A(\regs[8][10] ), .Y(n859) );
  MUX2X1 U1104 ( .B(n859), .A(n334), .S(n971), .Y(n1215) );
  INVX2 U1105 ( .A(\regs[11][10] ), .Y(n860) );
  MUX2X1 U1106 ( .B(n860), .A(n334), .S(n972), .Y(n1263) );
  INVX2 U1107 ( .A(\regs[10][10] ), .Y(n862) );
  MUX2X1 U1108 ( .B(n862), .A(n334), .S(n973), .Y(n1247) );
  AOI22X1 U1109 ( .A(n976), .B(\regs[9][10] ), .C(n975), .D(\regs[8][10] ), 
        .Y(n867) );
  AOI22X1 U1110 ( .A(n978), .B(\regs[11][10] ), .C(n977), .D(\regs[10][10] ), 
        .Y(n866) );
  INVX2 U1111 ( .A(\regs[13][10] ), .Y(n1429) );
  INVX2 U1112 ( .A(\regs[12][10] ), .Y(n1428) );
  OAI22X1 U1113 ( .A(n1429), .B(n544), .C(n1428), .D(n546), .Y(n864) );
  INVX2 U1114 ( .A(\regs[15][10] ), .Y(n1431) );
  INVX2 U1115 ( .A(\regs[14][10] ), .Y(n1430) );
  OAI22X1 U1116 ( .A(n1431), .B(n547), .C(n1430), .D(n549), .Y(n863) );
  NOR2X1 U1117 ( .A(n864), .B(n863), .Y(n865) );
  NAND3X1 U1118 ( .A(n867), .B(n866), .C(n865), .Y(n879) );
  AOI22X1 U1119 ( .A(\regs[7][10] ), .B(n514), .C(outreg_data[10]), .D(n884), 
        .Y(n877) );
  AOI22X1 U1136 ( .A(n406), .B(\regs[6][10] ), .C(n357), .D(\regs[1][10] ), 
        .Y(n876) );
  OAI22X1 U1153 ( .A(n870), .B(n869), .C(n868), .D(n1441), .Y(n874) );
  NOR2X1 U1170 ( .A(n873), .B(n874), .Y(n875) );
  NAND3X1 U1187 ( .A(n877), .B(n876), .C(n875), .Y(n878) );
  INVX2 U1188 ( .A(\regs[5][11] ), .Y(n1474) );
  INVX2 U1189 ( .A(\regs[2][11] ), .Y(n1465) );
  INVX2 U1190 ( .A(\regs[6][11] ), .Y(n1467) );
  INVX2 U1191 ( .A(\regs[7][11] ), .Y(n1476) );
  INVX2 U1192 ( .A(\regs[3][11] ), .Y(n1472) );
  INVX2 U1193 ( .A(\regs[9][11] ), .Y(n1461) );
  MUX2X1 U1194 ( .B(n1461), .A(n883), .S(n970), .Y(n1232) );
  INVX2 U1195 ( .A(\regs[8][11] ), .Y(n880) );
  MUX2X1 U1196 ( .B(n880), .A(n883), .S(n971), .Y(n1216) );
  INVX2 U1197 ( .A(\regs[11][11] ), .Y(n881) );
  MUX2X1 U1198 ( .B(n881), .A(n883), .S(n972), .Y(n1264) );
  INVX2 U1199 ( .A(\regs[10][11] ), .Y(n882) );
  MUX2X1 U1200 ( .B(n882), .A(n883), .S(n973), .Y(n1248) );
  INVX2 U1201 ( .A(\regs[4][11] ), .Y(n1466) );
  INVX2 U1202 ( .A(\regs[1][11] ), .Y(n1470) );
  AOI22X1 U1203 ( .A(n448), .B(\regs[5][11] ), .C(n422), .D(outreg_data[11]), 
        .Y(n899) );
  AOI22X1 U1204 ( .A(\regs[2][11] ), .B(n401), .C(n424), .D(\regs[6][11] ), 
        .Y(n898) );
  AOI22X1 U1205 ( .A(n548), .B(\regs[14][11] ), .C(n366), .D(\regs[15][11] ), 
        .Y(n886) );
  AOI22X1 U1206 ( .A(n545), .B(\regs[12][11] ), .C(n543), .D(\regs[13][11] ), 
        .Y(n885) );
  NAND2X1 U1207 ( .A(n886), .B(n885), .Y(n890) );
  AOI22X1 U1208 ( .A(n976), .B(\regs[9][11] ), .C(n975), .D(\regs[8][11] ), 
        .Y(n888) );
  AOI22X1 U1209 ( .A(n978), .B(\regs[11][11] ), .C(n977), .D(\regs[10][11] ), 
        .Y(n887) );
  NAND2X1 U1210 ( .A(n888), .B(n887), .Y(n889) );
  NOR2X1 U1211 ( .A(n890), .B(n889), .Y(n891) );
  OAI21X1 U1212 ( .A(n892), .B(n1472), .C(n891), .Y(n896) );
  AOI22X1 U1213 ( .A(n513), .B(\regs[4][11] ), .C(n893), .D(\regs[1][11] ), 
        .Y(n894) );
  OAI21X1 U1214 ( .A(n1476), .B(n539), .C(n894), .Y(n895) );
  NOR2X1 U1215 ( .A(n896), .B(n895), .Y(n897) );
  NAND3X1 U1216 ( .A(n898), .B(n899), .C(n897), .Y(r2_data[11]) );
  INVX2 U1217 ( .A(\regs[5][12] ), .Y(n900) );
  INVX2 U1218 ( .A(\regs[4][12] ), .Y(n901) );
  INVX2 U1219 ( .A(\regs[2][12] ), .Y(n902) );
  INVX2 U1220 ( .A(\regs[3][12] ), .Y(n903) );
  INVX2 U1221 ( .A(\regs[7][12] ), .Y(n912) );
  INVX2 U1222 ( .A(\regs[6][12] ), .Y(n913) );
  INVX2 U1223 ( .A(\regs[1][12] ), .Y(n911) );
  INVX2 U1224 ( .A(\regs[9][12] ), .Y(n1485) );
  MUX2X1 U1225 ( .B(n1485), .A(n330), .S(n970), .Y(n1233) );
  INVX2 U1226 ( .A(\regs[8][12] ), .Y(n1494) );
  MUX2X1 U1227 ( .B(n1494), .A(n330), .S(n971), .Y(n1217) );
  INVX2 U1228 ( .A(\regs[11][12] ), .Y(n1486) );
  MUX2X1 U1229 ( .B(n1486), .A(n330), .S(n972), .Y(n1265) );
  INVX2 U1230 ( .A(\regs[10][12] ), .Y(n1495) );
  MUX2X1 U1231 ( .B(n1495), .A(n330), .S(n973), .Y(n1249) );
  AOI22X1 U1232 ( .A(n976), .B(\regs[9][12] ), .C(n975), .D(\regs[8][12] ), 
        .Y(n909) );
  AOI22X1 U1233 ( .A(n978), .B(\regs[11][12] ), .C(n977), .D(\regs[10][12] ), 
        .Y(n908) );
  INVX2 U1234 ( .A(\regs[13][12] ), .Y(n1484) );
  INVX2 U1235 ( .A(\regs[12][12] ), .Y(n1493) );
  OAI22X1 U1236 ( .A(n1484), .B(n544), .C(n1493), .D(n546), .Y(n906) );
  INVX2 U1237 ( .A(\regs[15][12] ), .Y(n1483) );
  INVX2 U1238 ( .A(\regs[14][12] ), .Y(n1492) );
  OAI22X1 U1239 ( .A(n1483), .B(n547), .C(n1492), .D(n549), .Y(n905) );
  NOR2X1 U1240 ( .A(n906), .B(n905), .Y(n907) );
  NAND3X1 U1241 ( .A(n909), .B(n908), .C(n907), .Y(n920) );
  AOI22X1 U1242 ( .A(n448), .B(\regs[5][12] ), .C(n988), .D(\regs[4][12] ), 
        .Y(n918) );
  AOI22X1 U1243 ( .A(n398), .B(\regs[2][12] ), .C(n410), .D(\regs[3][12] ), 
        .Y(n917) );
  OAI22X1 U1244 ( .A(n911), .B(n430), .C(n910), .D(n358), .Y(n915) );
  OAI22X1 U1245 ( .A(n913), .B(n553), .C(n912), .D(n538), .Y(n914) );
  NOR2X1 U1246 ( .A(n915), .B(n914), .Y(n916) );
  NAND3X1 U1247 ( .A(n918), .B(n917), .C(n916), .Y(n919) );
  OR2X2 U1248 ( .A(n920), .B(n919), .Y(r2_data[12]) );
  INVX2 U1249 ( .A(\regs[5][13] ), .Y(n921) );
  INVX2 U1250 ( .A(\regs[4][13] ), .Y(n922) );
  INVX2 U1251 ( .A(\regs[2][13] ), .Y(n923) );
  INVX2 U1252 ( .A(\regs[3][13] ), .Y(n924) );
  INVX2 U1253 ( .A(\regs[7][13] ), .Y(n933) );
  INVX2 U1254 ( .A(\regs[6][13] ), .Y(n934) );
  INVX2 U1255 ( .A(\regs[1][13] ), .Y(n932) );
  INVX2 U1256 ( .A(\regs[9][13] ), .Y(n1505) );
  MUX2X1 U1257 ( .B(n1505), .A(n347), .S(n970), .Y(n1234) );
  INVX2 U1258 ( .A(\regs[8][13] ), .Y(n1514) );
  MUX2X1 U1259 ( .B(n1514), .A(n347), .S(n971), .Y(n1218) );
  INVX2 U1260 ( .A(\regs[11][13] ), .Y(n1506) );
  MUX2X1 U1261 ( .B(n1506), .A(n347), .S(n972), .Y(n1266) );
  INVX2 U1262 ( .A(\regs[10][13] ), .Y(n1515) );
  MUX2X1 U1263 ( .B(n1515), .A(n347), .S(n973), .Y(n1250) );
  AOI22X1 U1264 ( .A(n976), .B(\regs[9][13] ), .C(n975), .D(\regs[8][13] ), 
        .Y(n930) );
  AOI22X1 U1265 ( .A(n978), .B(\regs[11][13] ), .C(n977), .D(\regs[10][13] ), 
        .Y(n929) );
  INVX2 U1266 ( .A(\regs[13][13] ), .Y(n1504) );
  INVX2 U1267 ( .A(\regs[12][13] ), .Y(n1513) );
  OAI22X1 U1268 ( .A(n1504), .B(n544), .C(n1513), .D(n546), .Y(n927) );
  INVX2 U1269 ( .A(\regs[15][13] ), .Y(n1503) );
  INVX2 U1270 ( .A(\regs[14][13] ), .Y(n1512) );
  OAI22X1 U1271 ( .A(n1503), .B(n547), .C(n1512), .D(n549), .Y(n926) );
  NOR2X1 U1272 ( .A(n927), .B(n926), .Y(n928) );
  NAND3X1 U1273 ( .A(n930), .B(n929), .C(n928), .Y(n941) );
  AOI22X1 U1274 ( .A(n448), .B(\regs[5][13] ), .C(n988), .D(\regs[4][13] ), 
        .Y(n939) );
  AOI22X1 U1275 ( .A(n398), .B(\regs[2][13] ), .C(n410), .D(\regs[3][13] ), 
        .Y(n938) );
  OAI22X1 U1276 ( .A(n932), .B(n430), .C(n931), .D(n358), .Y(n936) );
  OAI22X1 U1277 ( .A(n934), .B(n553), .C(n321), .D(n933), .Y(n935) );
  NOR2X1 U1278 ( .A(n936), .B(n935), .Y(n937) );
  NAND3X1 U1279 ( .A(n939), .B(n938), .C(n937), .Y(n940) );
  OR2X2 U1280 ( .A(n941), .B(n940), .Y(r2_data[13]) );
  INVX2 U1281 ( .A(\regs[5][14] ), .Y(n942) );
  INVX2 U1282 ( .A(\regs[4][14] ), .Y(n943) );
  INVX2 U1283 ( .A(\regs[2][14] ), .Y(n944) );
  INVX2 U1284 ( .A(\regs[3][14] ), .Y(n945) );
  INVX2 U1285 ( .A(\regs[7][14] ), .Y(n954) );
  INVX2 U1286 ( .A(\regs[6][14] ), .Y(n955) );
  INVX2 U1287 ( .A(\regs[1][14] ), .Y(n953) );
  INVX2 U1288 ( .A(\regs[9][14] ), .Y(n1525) );
  MUX2X1 U1289 ( .B(n1525), .A(n336), .S(n970), .Y(n1235) );
  INVX2 U1290 ( .A(\regs[8][14] ), .Y(n1534) );
  MUX2X1 U1291 ( .B(n1534), .A(n336), .S(n971), .Y(n1219) );
  INVX2 U1292 ( .A(\regs[11][14] ), .Y(n1526) );
  MUX2X1 U1293 ( .B(n1526), .A(n336), .S(n972), .Y(n1267) );
  INVX2 U1294 ( .A(\regs[10][14] ), .Y(n1535) );
  MUX2X1 U1295 ( .B(n1535), .A(n336), .S(n973), .Y(n1251) );
  AOI22X1 U1296 ( .A(n976), .B(\regs[9][14] ), .C(n975), .D(\regs[8][14] ), 
        .Y(n951) );
  AOI22X1 U1297 ( .A(n978), .B(\regs[11][14] ), .C(n977), .D(\regs[10][14] ), 
        .Y(n950) );
  INVX2 U1298 ( .A(\regs[13][14] ), .Y(n1524) );
  INVX2 U1299 ( .A(\regs[12][14] ), .Y(n1533) );
  OAI22X1 U1301 ( .A(n1524), .B(n544), .C(n1533), .D(n546), .Y(n948) );
  INVX2 U1302 ( .A(\regs[15][14] ), .Y(n1523) );
  INVX2 U1303 ( .A(\regs[14][14] ), .Y(n1532) );
  OAI22X1 U1304 ( .A(n1523), .B(n547), .C(n1532), .D(n549), .Y(n947) );
  NOR2X1 U1305 ( .A(n948), .B(n947), .Y(n949) );
  NAND3X1 U1306 ( .A(n951), .B(n950), .C(n949), .Y(n962) );
  AOI22X1 U1307 ( .A(n448), .B(\regs[5][14] ), .C(n988), .D(\regs[4][14] ), 
        .Y(n960) );
  AOI22X1 U1308 ( .A(n416), .B(\regs[2][14] ), .C(n410), .D(\regs[3][14] ), 
        .Y(n959) );
  OAI22X1 U1309 ( .A(n953), .B(n430), .C(n952), .D(n358), .Y(n957) );
  OAI22X1 U1310 ( .A(n955), .B(n553), .C(n321), .D(n954), .Y(n956) );
  NOR2X1 U1311 ( .A(n957), .B(n956), .Y(n958) );
  NAND3X1 U1312 ( .A(n960), .B(n959), .C(n958), .Y(n961) );
  OR2X2 U1313 ( .A(n962), .B(n961), .Y(r2_data[14]) );
  INVX2 U1314 ( .A(\regs[5][15] ), .Y(n963) );
  MUX2X1 U1315 ( .B(n963), .A(n974), .S(n525), .Y(n1172) );
  INVX2 U1316 ( .A(\regs[4][15] ), .Y(n964) );
  MUX2X1 U1317 ( .B(n964), .A(n974), .S(n524), .Y(n1156) );
  INVX2 U1318 ( .A(\regs[2][15] ), .Y(n966) );
  MUX2X1 U1319 ( .B(n966), .A(n974), .S(n965), .Y(n465) );
  INVX2 U1320 ( .A(\regs[3][15] ), .Y(n968) );
  MUX2X1 U1321 ( .B(n968), .A(n974), .S(n967), .Y(n449) );
  INVX2 U1322 ( .A(\regs[7][15] ), .Y(n994) );
  MUX2X1 U1323 ( .B(n994), .A(n974), .S(n522), .Y(n1204) );
  INVX2 U1324 ( .A(\regs[6][15] ), .Y(n997) );
  MUX2X1 U1325 ( .B(n997), .A(n974), .S(n523), .Y(n1188) );
  INVX2 U1326 ( .A(\regs[1][15] ), .Y(n992) );
  MUX2X1 U1327 ( .B(n992), .A(n974), .S(n969), .Y(n481) );
  INVX2 U1328 ( .A(\regs[9][15] ), .Y(n1551) );
  MUX2X1 U1329 ( .B(n1551), .A(n335), .S(n970), .Y(n1236) );
  INVX2 U1330 ( .A(\regs[8][15] ), .Y(n1567) );
  MUX2X1 U1331 ( .B(n1567), .A(n335), .S(n971), .Y(n1220) );
  INVX2 U1332 ( .A(\regs[11][15] ), .Y(n1553) );
  MUX2X1 U1333 ( .B(n1553), .A(n974), .S(n972), .Y(n1268) );
  INVX2 U1334 ( .A(\regs[10][15] ), .Y(n1569) );
  MUX2X1 U1335 ( .B(n1569), .A(n335), .S(n973), .Y(n1252) );
  AOI22X1 U1336 ( .A(n976), .B(\regs[9][15] ), .C(n975), .D(\regs[8][15] ), 
        .Y(n987) );
  AOI22X1 U1337 ( .A(n978), .B(\regs[11][15] ), .C(n977), .D(\regs[10][15] ), 
        .Y(n986) );
  INVX2 U1338 ( .A(\regs[13][15] ), .Y(n1549) );
  INVX2 U1339 ( .A(\regs[12][15] ), .Y(n1565) );
  OAI22X1 U1340 ( .A(n1549), .B(n544), .C(n1565), .D(n546), .Y(n983) );
  INVX2 U1341 ( .A(\regs[15][15] ), .Y(n1547) );
  INVX2 U1342 ( .A(\regs[14][15] ), .Y(n1563) );
  OAI22X1 U1343 ( .A(n1547), .B(n547), .C(n1563), .D(n549), .Y(n982) );
  NOR2X1 U1344 ( .A(n983), .B(n982), .Y(n984) );
  NAND3X1 U1345 ( .A(n987), .B(n986), .C(n984), .Y(n1069) );
  AOI22X1 U1346 ( .A(n448), .B(\regs[5][15] ), .C(n988), .D(\regs[4][15] ), 
        .Y(n1035) );
  AOI22X1 U1347 ( .A(n432), .B(\regs[2][15] ), .C(n410), .D(\regs[3][15] ), 
        .Y(n1018) );
  OAI22X1 U1348 ( .A(n992), .B(n551), .C(n990), .D(n358), .Y(n1000) );
  OAI22X1 U1349 ( .A(n322), .B(n997), .C(n994), .D(n538), .Y(n998) );
  NOR2X1 U1350 ( .A(n1000), .B(n998), .Y(n1016) );
  NAND3X1 U1351 ( .A(n1035), .B(n1018), .C(n1016), .Y(n1053) );
  INVX2 U1352 ( .A(r1_sel[3]), .Y(n1071) );
  NAND2X1 U1353 ( .A(r1_sel[2]), .B(n1071), .Y(n1439) );
  NAND2X1 U1354 ( .A(n518), .B(n564), .Y(n1070) );
  NAND2X1 U1355 ( .A(n564), .B(n417), .Y(n1073) );
  AOI22X1 U1356 ( .A(\regs[7][0] ), .B(n1543), .C(\regs[3][0] ), .D(n1546), 
        .Y(n1095) );
  NAND2X1 U1357 ( .A(n405), .B(n1438), .Y(n1471) );
  NAND2X1 U1358 ( .A(n564), .B(n1361), .Y(n1074) );
  NAND3X1 U1359 ( .A(n565), .B(n985), .C(n1438), .Y(n1552) );
  NAND3X1 U1360 ( .A(n985), .B(n1438), .C(n393), .Y(n1568) );
  AOI22X1 U1361 ( .A(\regs[9][0] ), .B(n1318), .C(\regs[8][0] ), .D(n1459), 
        .Y(n1083) );
  NAND2X1 U1362 ( .A(n565), .B(n530), .Y(n1554) );
  NAND2X1 U1363 ( .A(n530), .B(n1315), .Y(n1570) );
  AOI22X1 U1364 ( .A(\regs[11][0] ), .B(n1458), .C(\regs[10][0] ), .D(n1453), 
        .Y(n1082) );
  NAND3X1 U1365 ( .A(n565), .B(n535), .C(n1438), .Y(n1550) );
  NAND3X1 U1366 ( .A(n535), .B(n1438), .C(n393), .Y(n1566) );
  OAI22X1 U1367 ( .A(n556), .B(n1076), .C(n558), .D(n1075), .Y(n1080) );
  NAND3X1 U1368 ( .A(n565), .B(n399), .C(n535), .Y(n1548) );
  NAND3X1 U1369 ( .A(n535), .B(n399), .C(n393), .Y(n1564) );
  OAI22X1 U1370 ( .A(n1548), .B(n1078), .C(n562), .D(n1077), .Y(n1079) );
  NOR2X1 U1371 ( .A(n1080), .B(n1079), .Y(n1081) );
  NAND3X1 U1372 ( .A(n1083), .B(n1082), .C(n1081), .Y(n1084) );
  AOI21X1 U1373 ( .A(\regs[1][0] ), .B(n385), .C(n1084), .Y(n1094) );
  NAND2X1 U1374 ( .A(n1361), .B(n1335), .Y(n1443) );
  OAI22X1 U1375 ( .A(n415), .B(n1086), .C(n419), .D(n1085), .Y(n1092) );
  NAND2X1 U1376 ( .A(n542), .B(n563), .Y(n1422) );
  NAND2X1 U1377 ( .A(n417), .B(n563), .Y(n1088) );
  AOI22X1 U1378 ( .A(\regs[4][0] ), .B(n1561), .C(\regs[2][0] ), .D(n1562), 
        .Y(n1089) );
  OAI21X1 U1379 ( .A(n412), .B(n1090), .C(n1089), .Y(n1091) );
  NOR2X1 U1380 ( .A(n1092), .B(n1091), .Y(n1093) );
  NAND3X1 U1381 ( .A(n1095), .B(n1094), .C(n1093), .Y(r1_data[0]) );
  NAND2X1 U1382 ( .A(n1375), .B(n1438), .Y(n1109) );
  OAI22X1 U1383 ( .A(n1471), .B(n1097), .C(n1473), .D(n1096), .Y(n1116) );
  AOI22X1 U1384 ( .A(\regs[9][1] ), .B(n1318), .C(\regs[8][1] ), .D(n1459), 
        .Y(n1106) );
  AOI22X1 U1385 ( .A(\regs[11][1] ), .B(n1458), .C(\regs[10][1] ), .D(n1453), 
        .Y(n1105) );
  INVX2 U1386 ( .A(\regs[13][1] ), .Y(n1099) );
  INVX2 U1387 ( .A(\regs[12][1] ), .Y(n1098) );
  OAI22X1 U1388 ( .A(n556), .B(n1099), .C(n1566), .D(n1098), .Y(n1103) );
  INVX2 U1389 ( .A(\regs[15][1] ), .Y(n1101) );
  INVX2 U1390 ( .A(\regs[14][1] ), .Y(n1100) );
  OAI22X1 U1391 ( .A(n560), .B(n1101), .C(n1564), .D(n1100), .Y(n1102) );
  NOR2X1 U1392 ( .A(n1103), .B(n1102), .Y(n1104) );
  NAND3X1 U1393 ( .A(n1106), .B(n1105), .C(n1104), .Y(n1110) );
  INVX2 U1394 ( .A(n1110), .Y(n1108) );
  NAND2X1 U1395 ( .A(n537), .B(n1438), .Y(n1119) );
  INVX2 U1396 ( .A(n1119), .Y(n1132) );
  AOI22X1 U1397 ( .A(\regs[6][1] ), .B(n518), .C(\regs[4][1] ), .D(n1132), .Y(
        n1107) );
  NAND3X1 U1398 ( .A(n1108), .B(n391), .C(n1107), .Y(n1115) );
  AOI22X1 U1399 ( .A(\regs[3][1] ), .B(n433), .C(\regs[1][1] ), .D(n407), .Y(
        n1113) );
  AOI22X1 U1400 ( .A(\regs[7][1] ), .B(n518), .C(n1132), .D(\regs[5][1] ), .Y(
        n1112) );
  NOR2X1 U1401 ( .A(n1335), .B(n1110), .Y(n1111) );
  NAND3X1 U1402 ( .A(n1113), .B(n1112), .C(n1111), .Y(n1114) );
  OAI21X1 U1403 ( .A(n1116), .B(n1115), .C(n1114), .Y(n1117) );
  INVX2 U1404 ( .A(n1117), .Y(r1_data[1]) );
  OAI22X1 U1405 ( .A(n1477), .B(n1120), .C(n384), .D(n1118), .Y(n1139) );
  AOI22X1 U1406 ( .A(\regs[9][2] ), .B(n1318), .C(\regs[8][2] ), .D(n1459), 
        .Y(n1129) );
  AOI22X1 U1407 ( .A(\regs[11][2] ), .B(n1458), .C(\regs[10][2] ), .D(n1453), 
        .Y(n1128) );
  OAI22X1 U1408 ( .A(n556), .B(n1122), .C(n558), .D(n1121), .Y(n1126) );
  OAI22X1 U1409 ( .A(n1548), .B(n1124), .C(n562), .D(n1123), .Y(n1125) );
  NOR2X1 U1410 ( .A(n1126), .B(n1125), .Y(n1127) );
  NAND3X1 U1411 ( .A(n1129), .B(n1128), .C(n1127), .Y(n1133) );
  INVX2 U1412 ( .A(n1133), .Y(n1131) );
  AOI22X1 U1413 ( .A(\regs[1][2] ), .B(n361), .C(\regs[3][2] ), .D(n433), .Y(
        n1130) );
  NAND3X1 U1414 ( .A(n1131), .B(n565), .C(n1130), .Y(n1138) );
  AOI22X1 U1415 ( .A(n361), .B(outreg_data[2]), .C(n433), .D(\regs[2][2] ), 
        .Y(n1136) );
  AOI22X1 U1416 ( .A(n1132), .B(\regs[4][2] ), .C(\regs[6][2] ), .D(n542), .Y(
        n1135) );
  NAND3X1 U1417 ( .A(n1134), .B(n1136), .C(n1135), .Y(n1137) );
  OAI21X1 U1418 ( .A(n1139), .B(n1138), .C(n1137), .Y(n1269) );
  INVX2 U1419 ( .A(n1269), .Y(r1_data[2]) );
  OAI22X1 U1420 ( .A(n1477), .B(n1271), .C(n447), .D(n1270), .Y(n1275) );
  OAI22X1 U1421 ( .A(n1473), .B(n1273), .C(n411), .D(n1272), .Y(n1274) );
  NOR2X1 U1422 ( .A(n1275), .B(n1274), .Y(n1295) );
  AOI22X1 U1423 ( .A(\regs[9][3] ), .B(n1318), .C(\regs[8][3] ), .D(n1459), 
        .Y(n1284) );
  AOI22X1 U1424 ( .A(\regs[11][3] ), .B(n1458), .C(\regs[10][3] ), .D(n1453), 
        .Y(n1283) );
  OAI22X1 U1425 ( .A(n1550), .B(n1277), .C(n1566), .D(n1276), .Y(n1281) );
  OAI22X1 U1426 ( .A(n560), .B(n1279), .C(n1564), .D(n1278), .Y(n1280) );
  NOR2X1 U1427 ( .A(n1281), .B(n1280), .Y(n1282) );
  NAND3X1 U1428 ( .A(n1284), .B(n1283), .C(n1282), .Y(n1291) );
  NOR2X1 U1429 ( .A(n391), .B(n1291), .Y(n1294) );
  OAI22X1 U1430 ( .A(n1477), .B(n1286), .C(n447), .D(n1285), .Y(n1290) );
  OAI22X1 U1431 ( .A(n1473), .B(n1288), .C(n1471), .D(n1287), .Y(n1289) );
  NOR2X1 U1432 ( .A(n1290), .B(n1289), .Y(n1293) );
  NOR2X1 U1433 ( .A(n565), .B(n1291), .Y(n1292) );
  AOI22X1 U1434 ( .A(n1295), .B(n1294), .C(n1293), .D(n1292), .Y(r1_data[3])
         );
  AOI22X1 U1435 ( .A(\regs[7][4] ), .B(n1543), .C(\regs[3][4] ), .D(n1546), 
        .Y(n1314) );
  AOI22X1 U1436 ( .A(\regs[9][4] ), .B(n1318), .C(\regs[8][4] ), .D(n1459), 
        .Y(n1304) );
  AOI22X1 U1437 ( .A(\regs[11][4] ), .B(n1458), .C(\regs[10][4] ), .D(n1453), 
        .Y(n1303) );
  OAI22X1 U1438 ( .A(n556), .B(n1297), .C(n558), .D(n1296), .Y(n1301) );
  OAI22X1 U1439 ( .A(n1548), .B(n1299), .C(n562), .D(n1298), .Y(n1300) );
  NOR2X1 U1440 ( .A(n1301), .B(n1300), .Y(n1302) );
  NAND3X1 U1441 ( .A(n1304), .B(n1303), .C(n1302), .Y(n1305) );
  AOI21X1 U1442 ( .A(n1545), .B(\regs[1][4] ), .C(n1305), .Y(n1313) );
  OAI22X1 U1443 ( .A(n415), .B(n1307), .C(n419), .D(n1306), .Y(n1311) );
  AOI22X1 U1444 ( .A(\regs[4][4] ), .B(n1561), .C(\regs[2][4] ), .D(n1562), 
        .Y(n1308) );
  NOR2X1 U1445 ( .A(n1310), .B(n1311), .Y(n1312) );
  AOI22X1 U1446 ( .A(n417), .B(\regs[3][5] ), .C(\regs[7][5] ), .D(n518), .Y(
        n1317) );
  NAND2X1 U1447 ( .A(\regs[1][5] ), .B(n407), .Y(n1316) );
  AOI21X1 U1448 ( .A(n1317), .B(n1316), .C(n1315), .Y(n1332) );
  INVX2 U1449 ( .A(n1552), .Y(n1318) );
  AOI22X1 U1450 ( .A(\regs[9][5] ), .B(n1318), .C(\regs[8][5] ), .D(n1459), 
        .Y(n1320) );
  AOI22X1 U1451 ( .A(\regs[11][5] ), .B(n1458), .C(\regs[10][5] ), .D(n1453), 
        .Y(n1319) );
  NAND2X1 U1452 ( .A(n1320), .B(n1319), .Y(n1331) );
  NAND3X1 U1453 ( .A(outreg_data[5]), .B(n361), .C(n1315), .Y(n1329) );
  NAND3X1 U1454 ( .A(\regs[5][5] ), .B(n446), .C(n565), .Y(n1328) );
  OAI22X1 U1455 ( .A(n1550), .B(n1322), .C(n1566), .D(n1321), .Y(n1326) );
  OAI22X1 U1456 ( .A(n560), .B(n1324), .C(n1564), .D(n1323), .Y(n1325) );
  NOR2X1 U1457 ( .A(n1326), .B(n1325), .Y(n1327) );
  NAND3X1 U1458 ( .A(n1329), .B(n1328), .C(n1327), .Y(n1330) );
  NOR3X1 U1459 ( .A(n1331), .B(n1332), .C(n1330), .Y(n1339) );
  OAI22X1 U1460 ( .A(n1473), .B(n1334), .C(n1477), .D(n1333), .Y(n1337) );
  AND2X2 U1461 ( .A(\regs[4][5] ), .B(n446), .Y(n1336) );
  OAI21X1 U1462 ( .A(n1337), .B(n1336), .C(n1315), .Y(n1338) );
  NAND2X1 U1463 ( .A(n1339), .B(n1338), .Y(r1_data[5]) );
  OAI22X1 U1464 ( .A(n447), .B(n1341), .C(n1477), .D(n1340), .Y(n1359) );
  AOI22X1 U1465 ( .A(\regs[9][6] ), .B(n1318), .C(\regs[8][6] ), .D(n1459), 
        .Y(n1350) );
  AOI22X1 U1466 ( .A(\regs[11][6] ), .B(n1458), .C(\regs[10][6] ), .D(n1453), 
        .Y(n1349) );
  INVX2 U1467 ( .A(\regs[13][6] ), .Y(n1343) );
  INVX2 U1468 ( .A(\regs[12][6] ), .Y(n1342) );
  OAI22X1 U1469 ( .A(n556), .B(n1343), .C(n558), .D(n1342), .Y(n1347) );
  INVX2 U1470 ( .A(\regs[15][6] ), .Y(n1345) );
  INVX2 U1471 ( .A(\regs[14][6] ), .Y(n1344) );
  OAI22X1 U1472 ( .A(n1548), .B(n1345), .C(n562), .D(n1344), .Y(n1346) );
  NOR2X1 U1473 ( .A(n1347), .B(n1346), .Y(n1348) );
  NAND3X1 U1474 ( .A(n1350), .B(n1349), .C(n1348), .Y(n1353) );
  INVX2 U1475 ( .A(n1353), .Y(n1352) );
  AOI22X1 U1476 ( .A(outreg_data[6]), .B(n407), .C(\regs[2][6] ), .D(n433), 
        .Y(n1351) );
  NAND3X1 U1477 ( .A(n1352), .B(n391), .C(n1351), .Y(n1358) );
  AOI22X1 U1478 ( .A(\regs[1][6] ), .B(n361), .C(n433), .D(\regs[3][6] ), .Y(
        n1356) );
  AOI22X1 U1479 ( .A(\regs[5][6] ), .B(n446), .C(\regs[7][6] ), .D(n404), .Y(
        n1355) );
  NOR2X1 U1480 ( .A(n563), .B(n1353), .Y(n1354) );
  NAND3X1 U1481 ( .A(n1356), .B(n1354), .C(n1355), .Y(n1357) );
  OAI21X1 U1482 ( .A(n1359), .B(n1358), .C(n1357), .Y(n1360) );
  INVX2 U1483 ( .A(n1360), .Y(r1_data[6]) );
  NAND2X1 U1484 ( .A(\regs[7][7] ), .B(n1543), .Y(n1387) );
  NAND3X1 U1485 ( .A(n361), .B(n391), .C(outreg_data[7]), .Y(n1362) );
  INVX2 U1486 ( .A(n1362), .Y(n1384) );
  NAND3X1 U1487 ( .A(n446), .B(n565), .C(\regs[5][7] ), .Y(n1363) );
  INVX2 U1488 ( .A(n1363), .Y(n1383) );
  NAND2X1 U1489 ( .A(\regs[11][7] ), .B(n1458), .Y(n1365) );
  NAND2X1 U1490 ( .A(\regs[10][7] ), .B(n1453), .Y(n1364) );
  NAND2X1 U1491 ( .A(n1365), .B(n1364), .Y(n1372) );
  OAI22X1 U1492 ( .A(n1550), .B(n1367), .C(n1566), .D(n1366), .Y(n1371) );
  OAI22X1 U1493 ( .A(n560), .B(n1369), .C(n1564), .D(n1368), .Y(n1370) );
  NOR3X1 U1494 ( .A(n1372), .B(n1371), .C(n1370), .Y(n1381) );
  AOI22X1 U1495 ( .A(\regs[8][7] ), .B(n1459), .C(\regs[9][7] ), .D(n1318), 
        .Y(n1380) );
  NAND2X1 U1496 ( .A(\regs[6][7] ), .B(r1_sel[1]), .Y(n1374) );
  NAND2X1 U1497 ( .A(\regs[4][7] ), .B(n1438), .Y(n1373) );
  AOI21X1 U1498 ( .A(n1374), .B(n1373), .C(n439), .Y(n1378) );
  NAND3X1 U1499 ( .A(n390), .B(n405), .C(\regs[2][7] ), .Y(n1376) );
  INVX2 U1500 ( .A(n1376), .Y(n1377) );
  OAI21X1 U1501 ( .A(n1378), .B(n1377), .C(n391), .Y(n1379) );
  NAND3X1 U1502 ( .A(n1381), .B(n1380), .C(n1379), .Y(n1382) );
  NOR3X1 U1503 ( .A(n1384), .B(n1383), .C(n1382), .Y(n1386) );
  AOI22X1 U1504 ( .A(n1545), .B(\regs[1][7] ), .C(n1546), .D(\regs[3][7] ), 
        .Y(n1385) );
  NAND3X1 U1505 ( .A(n1385), .B(n1387), .C(n1386), .Y(r1_data[7]) );
  AOI22X1 U1506 ( .A(\regs[5][8] ), .B(n1544), .C(\regs[7][8] ), .D(n1543), 
        .Y(n1396) );
  AOI22X1 U1507 ( .A(n1546), .B(\regs[3][8] ), .C(n1545), .D(\regs[1][8] ), 
        .Y(n1395) );
  OAI22X1 U1508 ( .A(n556), .B(n1389), .C(n560), .D(n1388), .Y(n1393) );
  OAI22X1 U1509 ( .A(n1554), .B(n1391), .C(n1552), .D(n1390), .Y(n1392) );
  NOR2X1 U1510 ( .A(n1393), .B(n1392), .Y(n1394) );
  NAND3X1 U1511 ( .A(n1396), .B(n1395), .C(n1394), .Y(n1407) );
  AOI22X1 U1512 ( .A(\regs[4][8] ), .B(n1561), .C(\regs[6][8] ), .D(n1560), 
        .Y(n1405) );
  AOI22X1 U1513 ( .A(\regs[2][8] ), .B(n1562), .C(outreg_data[8]), .D(n541), 
        .Y(n1404) );
  OAI22X1 U1514 ( .A(n558), .B(n1398), .C(n562), .D(n1397), .Y(n1402) );
  OAI22X1 U1515 ( .A(n1570), .B(n1400), .C(n1568), .D(n1399), .Y(n1401) );
  NOR2X1 U1516 ( .A(n1402), .B(n1401), .Y(n1403) );
  NAND3X1 U1517 ( .A(n1405), .B(n1404), .C(n1403), .Y(n1406) );
  OR2X2 U1518 ( .A(n1406), .B(n1407), .Y(r1_data[8]) );
  AOI22X1 U1519 ( .A(\regs[7][9] ), .B(n1543), .C(\regs[3][9] ), .D(n1546), 
        .Y(n1427) );
  AOI22X1 U1520 ( .A(\regs[9][9] ), .B(n1318), .C(\regs[8][9] ), .D(n1459), 
        .Y(n1416) );
  AOI22X1 U1521 ( .A(\regs[11][9] ), .B(n1458), .C(\regs[10][9] ), .D(n1453), 
        .Y(n1415) );
  OAI22X1 U1522 ( .A(n1550), .B(n1409), .C(n558), .D(n1408), .Y(n1413) );
  OAI22X1 U1523 ( .A(n1548), .B(n1411), .C(n1564), .D(n1410), .Y(n1412) );
  NOR2X1 U1524 ( .A(n1413), .B(n1412), .Y(n1414) );
  NAND3X1 U1525 ( .A(n1416), .B(n1415), .C(n1414), .Y(n1417) );
  AOI21X1 U1526 ( .A(\regs[1][9] ), .B(n1545), .C(n1417), .Y(n1426) );
  OAI22X1 U1527 ( .A(n415), .B(n1419), .C(n377), .D(n1418), .Y(n1424) );
  AOI22X1 U1528 ( .A(\regs[4][9] ), .B(n1561), .C(\regs[2][9] ), .D(n1562), 
        .Y(n1420) );
  NOR2X1 U1529 ( .A(n1423), .B(n1424), .Y(n1425) );
  AOI22X1 U1530 ( .A(\regs[7][10] ), .B(n1543), .C(\regs[3][10] ), .D(n1546), 
        .Y(n1450) );
  AOI22X1 U1531 ( .A(\regs[9][10] ), .B(n1318), .C(\regs[8][10] ), .D(n1459), 
        .Y(n1436) );
  AOI22X1 U1532 ( .A(\regs[11][10] ), .B(n1458), .C(\regs[10][10] ), .D(n1453), 
        .Y(n1435) );
  OAI22X1 U1533 ( .A(n556), .B(n1429), .C(n1566), .D(n1428), .Y(n1433) );
  OAI22X1 U1534 ( .A(n560), .B(n1431), .C(n562), .D(n1430), .Y(n1432) );
  NOR2X1 U1535 ( .A(n1433), .B(n1432), .Y(n1434) );
  NAND3X1 U1536 ( .A(n1436), .B(n1435), .C(n1434), .Y(n1437) );
  AOI21X1 U1537 ( .A(n1545), .B(\regs[1][10] ), .C(n1437), .Y(n1449) );
  AOI22X1 U1538 ( .A(\regs[6][10] ), .B(n390), .C(\regs[4][10] ), .D(n1438), 
        .Y(n1440) );
  OAI22X1 U1539 ( .A(n1473), .B(n1441), .C(n1440), .D(n439), .Y(n1447) );
  OAI22X1 U1540 ( .A(n1445), .B(n1444), .C(n1443), .D(n1442), .Y(n1446) );
  AOI21X1 U1541 ( .A(n1447), .B(n393), .C(n1446), .Y(n1448) );
  NAND3X1 U1542 ( .A(n1450), .B(n1449), .C(n1448), .Y(r1_data[10]) );
  INVX2 U1543 ( .A(\regs[13][11] ), .Y(n1452) );
  INVX2 U1544 ( .A(\regs[12][11] ), .Y(n1451) );
  OAI22X1 U1545 ( .A(n1550), .B(n1452), .C(n558), .D(n1451), .Y(n1457) );
  INVX2 U1546 ( .A(\regs[15][11] ), .Y(n1455) );
  AOI22X1 U1547 ( .A(\regs[10][11] ), .B(n1453), .C(\regs[14][11] ), .D(n561), 
        .Y(n1454) );
  OAI21X1 U1548 ( .A(n560), .B(n1455), .C(n1454), .Y(n1456) );
  OR2X2 U1549 ( .A(n1457), .B(n1456), .Y(n1463) );
  AOI22X1 U1550 ( .A(\regs[8][11] ), .B(n1459), .C(\regs[11][11] ), .D(n1458), 
        .Y(n1460) );
  OAI21X1 U1551 ( .A(n1552), .B(n1461), .C(n1460), .Y(n1462) );
  NOR2X1 U1552 ( .A(n1463), .B(n1462), .Y(n1482) );
  OAI22X1 U1553 ( .A(n1473), .B(n1465), .C(n1464), .D(n1471), .Y(n1469) );
  OAI22X1 U1554 ( .A(n1477), .B(n1467), .C(n447), .D(n1466), .Y(n1468) );
  OAI21X1 U1555 ( .A(n1468), .B(n1469), .C(n393), .Y(n1481) );
  OAI22X1 U1556 ( .A(n1473), .B(n1472), .C(n1471), .D(n1470), .Y(n1479) );
  OAI22X1 U1557 ( .A(n1477), .B(n1476), .C(n447), .D(n1474), .Y(n1478) );
  OAI21X1 U1558 ( .A(n1479), .B(n1478), .C(n565), .Y(n1480) );
  NAND3X1 U1559 ( .A(n1482), .B(n1481), .C(n1480), .Y(r1_data[11]) );
  AOI22X1 U1560 ( .A(\regs[5][12] ), .B(n1544), .C(\regs[7][12] ), .D(n388), 
        .Y(n1491) );
  AOI22X1 U1561 ( .A(n1546), .B(\regs[3][12] ), .C(\regs[1][12] ), .D(n385), 
        .Y(n1490) );
  OAI22X1 U1562 ( .A(n556), .B(n1484), .C(n1548), .D(n1483), .Y(n1488) );
  OAI22X1 U1563 ( .A(n1554), .B(n1486), .C(n1552), .D(n1485), .Y(n1487) );
  NOR2X1 U1564 ( .A(n1488), .B(n1487), .Y(n1489) );
  NAND3X1 U1565 ( .A(n1491), .B(n1489), .C(n1490), .Y(n1502) );
  AOI22X1 U1566 ( .A(\regs[4][12] ), .B(n1561), .C(\regs[6][12] ), .D(n1560), 
        .Y(n1500) );
  AOI22X1 U1567 ( .A(\regs[2][12] ), .B(n1562), .C(outreg_data[12]), .D(n541), 
        .Y(n1499) );
  OAI22X1 U1568 ( .A(n558), .B(n1493), .C(n1564), .D(n1492), .Y(n1497) );
  OAI22X1 U1569 ( .A(n1570), .B(n1495), .C(n1568), .D(n1494), .Y(n1496) );
  NOR2X1 U1570 ( .A(n1497), .B(n1496), .Y(n1498) );
  NAND3X1 U1571 ( .A(n1500), .B(n1499), .C(n1498), .Y(n1501) );
  OR2X2 U1572 ( .A(n1502), .B(n1501), .Y(r1_data[12]) );
  AOI22X1 U1573 ( .A(\regs[5][13] ), .B(n1544), .C(\regs[7][13] ), .D(n1543), 
        .Y(n1511) );
  AOI22X1 U1574 ( .A(n1546), .B(\regs[3][13] ), .C(n1545), .D(\regs[1][13] ), 
        .Y(n1510) );
  OAI22X1 U1575 ( .A(n1550), .B(n1504), .C(n560), .D(n1503), .Y(n1508) );
  OAI22X1 U1576 ( .A(n1554), .B(n1506), .C(n1552), .D(n1505), .Y(n1507) );
  NOR2X1 U1577 ( .A(n1508), .B(n1507), .Y(n1509) );
  NAND3X1 U1578 ( .A(n1511), .B(n1510), .C(n1509), .Y(n1522) );
  AOI22X1 U1579 ( .A(\regs[4][13] ), .B(n1561), .C(\regs[6][13] ), .D(n420), 
        .Y(n1520) );
  AOI22X1 U1580 ( .A(\regs[2][13] ), .B(n1562), .C(outreg_data[13]), .D(n541), 
        .Y(n1519) );
  OAI22X1 U1581 ( .A(n1566), .B(n1513), .C(n562), .D(n1512), .Y(n1517) );
  OAI22X1 U1582 ( .A(n1570), .B(n1515), .C(n1568), .D(n1514), .Y(n1516) );
  NOR2X1 U1583 ( .A(n1517), .B(n1516), .Y(n1518) );
  NAND3X1 U1584 ( .A(n1518), .B(n1519), .C(n1520), .Y(n1521) );
  OR2X2 U1585 ( .A(n1521), .B(n1522), .Y(r1_data[13]) );
  AOI22X1 U1586 ( .A(\regs[5][14] ), .B(n1544), .C(\regs[7][14] ), .D(n1543), 
        .Y(n1531) );
  AOI22X1 U1587 ( .A(\regs[3][14] ), .B(n1546), .C(\regs[1][14] ), .D(n385), 
        .Y(n1530) );
  OAI22X1 U1588 ( .A(n556), .B(n1524), .C(n1548), .D(n1523), .Y(n1528) );
  OAI22X1 U1589 ( .A(n1554), .B(n1526), .C(n1552), .D(n1525), .Y(n1527) );
  NOR2X1 U1590 ( .A(n1528), .B(n1527), .Y(n1529) );
  NAND3X1 U1591 ( .A(n1530), .B(n1531), .C(n1529), .Y(n1542) );
  AOI22X1 U1592 ( .A(\regs[4][14] ), .B(n1561), .C(\regs[6][14] ), .D(n1560), 
        .Y(n1540) );
  AOI22X1 U1593 ( .A(n1562), .B(\regs[2][14] ), .C(outreg_data[14]), .D(n541), 
        .Y(n1539) );
  OAI22X1 U1594 ( .A(n558), .B(n1533), .C(n1564), .D(n1532), .Y(n1537) );
  OAI22X1 U1595 ( .A(n1570), .B(n1535), .C(n1568), .D(n1534), .Y(n1536) );
  NOR2X1 U1596 ( .A(n1537), .B(n1536), .Y(n1538) );
  NAND3X1 U1597 ( .A(n1539), .B(n1540), .C(n1538), .Y(n1541) );
  OR2X2 U1598 ( .A(n1542), .B(n1541), .Y(r1_data[14]) );
  AOI22X1 U1599 ( .A(\regs[5][15] ), .B(n1544), .C(\regs[7][15] ), .D(n1543), 
        .Y(n1559) );
  AOI22X1 U1600 ( .A(\regs[3][15] ), .B(n1546), .C(n1545), .D(\regs[1][15] ), 
        .Y(n1558) );
  OAI22X1 U1601 ( .A(n1550), .B(n1549), .C(n560), .D(n1547), .Y(n1556) );
  OAI22X1 U1602 ( .A(n1554), .B(n1553), .C(n1552), .D(n1551), .Y(n1555) );
  NOR2X1 U1603 ( .A(n1556), .B(n1555), .Y(n1557) );
  NAND3X1 U1604 ( .A(n1559), .B(n1558), .C(n1557), .Y(n1577) );
  AOI22X1 U1605 ( .A(\regs[4][15] ), .B(n1561), .C(\regs[6][15] ), .D(n1560), 
        .Y(n1575) );
  AOI22X1 U1606 ( .A(\regs[2][15] ), .B(n1562), .C(outreg_data[15]), .D(n541), 
        .Y(n1574) );
  OAI22X1 U1607 ( .A(n1566), .B(n1565), .C(n562), .D(n1563), .Y(n1572) );
  OAI22X1 U1608 ( .A(n1570), .B(n1569), .C(n1568), .D(n1567), .Y(n1571) );
  NOR2X1 U1609 ( .A(n1572), .B(n1571), .Y(n1573) );
  NAND3X1 U1610 ( .A(n1575), .B(n1574), .C(n1573), .Y(n1576) );
  OR2X2 U1611 ( .A(n1577), .B(n1576), .Y(r1_data[15]) );
endmodule


module scalable_cla_block_CLA_BLK_SIZE_BITS4_3 ( A, B, Cin, S, PG, GG );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  INVX2 U1 ( .A(A[1]), .Y(n37) );
  INVX4 U2 ( .A(A[3]), .Y(n35) );
  INVX1 U3 ( .A(n6), .Y(n3) );
  OR2X2 U4 ( .A(n3), .B(A[2]), .Y(n12) );
  NOR2X1 U5 ( .A(A[1]), .B(B[1]), .Y(n20) );
  INVX1 U6 ( .A(A[1]), .Y(n17) );
  INVX1 U7 ( .A(B[1]), .Y(n22) );
  INVX2 U8 ( .A(B[3]), .Y(n1) );
  INVX1 U9 ( .A(B[3]), .Y(n34) );
  BUFX2 U10 ( .A(B[0]), .Y(n2) );
  INVX2 U11 ( .A(B[2]), .Y(n6) );
  INVX1 U12 ( .A(n11), .Y(n4) );
  INVX1 U13 ( .A(n35), .Y(n8) );
  INVX1 U14 ( .A(n1), .Y(n11) );
  NAND2X1 U15 ( .A(n6), .B(n5), .Y(n44) );
  INVX1 U16 ( .A(A[2]), .Y(n5) );
  INVX1 U17 ( .A(n16), .Y(n7) );
  INVX1 U18 ( .A(n40), .Y(n9) );
  BUFX2 U19 ( .A(n44), .Y(n10) );
  AND2X2 U20 ( .A(A[2]), .B(B[2]), .Y(n13) );
  AND2X1 U21 ( .A(n44), .B(B[0]), .Y(n27) );
  INVX1 U22 ( .A(n13), .Y(n40) );
  INVX1 U23 ( .A(n17), .Y(n14) );
  BUFX2 U24 ( .A(A[0]), .Y(n15) );
  BUFX2 U25 ( .A(n18), .Y(n16) );
  INVX1 U26 ( .A(n22), .Y(n18) );
  BUFX2 U27 ( .A(n15), .Y(n19) );
  XNOR2X1 U28 ( .A(Cin), .B(n21), .Y(S[0]) );
  XNOR2X1 U29 ( .A(n15), .B(n2), .Y(n21) );
  INVX1 U30 ( .A(B[1]), .Y(n36) );
  OAI21X1 U31 ( .A(A[3]), .B(B[3]), .C(n13), .Y(n24) );
  NAND2X1 U32 ( .A(B[3]), .B(A[3]), .Y(n23) );
  AND2X2 U33 ( .A(n24), .B(n23), .Y(n31) );
  NOR2X1 U34 ( .A(n37), .B(n36), .Y(n26) );
  NAND2X1 U35 ( .A(n35), .B(n34), .Y(n25) );
  NAND3X1 U36 ( .A(n26), .B(n25), .C(n12), .Y(n30) );
  NAND2X1 U37 ( .A(n37), .B(n7), .Y(n32) );
  AOI21X1 U38 ( .A(n35), .B(n1), .C(n20), .Y(n28) );
  NAND3X1 U39 ( .A(A[0]), .B(n27), .C(n28), .Y(n29) );
  NAND3X1 U40 ( .A(n31), .B(n29), .C(n30), .Y(GG) );
  NAND2X1 U41 ( .A(n32), .B(n10), .Y(n33) );
  AOI21X1 U42 ( .A(n35), .B(n4), .C(n33), .Y(PG) );
  OAI21X1 U43 ( .A(n19), .B(n2), .C(Cin), .Y(n47) );
  NAND2X1 U44 ( .A(A[0]), .B(B[0]), .Y(n46) );
  NAND2X1 U45 ( .A(n47), .B(n46), .Y(n38) );
  FAX1 U46 ( .A(n16), .B(n38), .C(n14), .YS(S[1]) );
  NAND2X1 U47 ( .A(n18), .B(n14), .Y(n45) );
  INVX2 U48 ( .A(n45), .Y(n39) );
  NAND2X1 U49 ( .A(n22), .B(n37), .Y(n43) );
  OAI21X1 U50 ( .A(n39), .B(n38), .C(n43), .Y(n42) );
  NAND2X1 U51 ( .A(n12), .B(n40), .Y(n41) );
  XOR2X1 U52 ( .A(n42), .B(n41), .Y(S[2]) );
  AND2X2 U53 ( .A(n43), .B(n10), .Y(n49) );
  NAND3X1 U54 ( .A(n47), .B(n46), .C(n45), .Y(n48) );
  AOI21X1 U55 ( .A(n49), .B(n48), .C(n9), .Y(n51) );
  XOR2X1 U56 ( .A(n11), .B(n8), .Y(n50) );
  XNOR2X1 U57 ( .A(n51), .B(n50), .Y(S[3]) );
endmodule


module scalable_cla_block_CLA_BLK_SIZE_BITS4_0 ( A, B, Cin, S, PG, GG );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output PG, GG;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66;

  AND2X2 U1 ( .A(n16), .B(n21), .Y(PG) );
  AND2X2 U2 ( .A(n11), .B(n32), .Y(n2) );
  AND2X2 U3 ( .A(n44), .B(n60), .Y(n3) );
  NAND2X1 U4 ( .A(n8), .B(n3), .Y(n45) );
  INVX4 U5 ( .A(B[3]), .Y(n48) );
  INVX1 U6 ( .A(A[3]), .Y(n25) );
  AND2X1 U7 ( .A(n63), .B(n62), .Y(n4) );
  NOR2X1 U8 ( .A(n4), .B(n61), .Y(n64) );
  AND2X2 U9 ( .A(n15), .B(n60), .Y(n6) );
  INVX2 U10 ( .A(n38), .Y(n60) );
  AND2X2 U11 ( .A(n27), .B(n10), .Y(n5) );
  AND2X2 U12 ( .A(n51), .B(n11), .Y(n7) );
  INVX1 U13 ( .A(Cin), .Y(n8) );
  INVX1 U14 ( .A(Cin), .Y(n14) );
  NAND2X1 U15 ( .A(n26), .B(n19), .Y(n9) );
  INVX2 U16 ( .A(B[1]), .Y(n26) );
  AND2X2 U17 ( .A(n54), .B(n53), .Y(n16) );
  BUFX2 U18 ( .A(n37), .Y(n10) );
  NAND2X1 U19 ( .A(n29), .B(n28), .Y(n11) );
  BUFX2 U20 ( .A(A[0]), .Y(n12) );
  INVX1 U21 ( .A(n10), .Y(n31) );
  NAND2X1 U22 ( .A(n37), .B(n36), .Y(n13) );
  INVX1 U23 ( .A(Cin), .Y(n49) );
  INVX1 U24 ( .A(n11), .Y(n30) );
  INVX1 U25 ( .A(n56), .Y(n57) );
  NAND2X1 U26 ( .A(Cin), .B(n7), .Y(n65) );
  INVX1 U27 ( .A(n59), .Y(n51) );
  INVX1 U28 ( .A(A[1]), .Y(n19) );
  INVX1 U29 ( .A(n53), .Y(n20) );
  INVX1 U30 ( .A(A[0]), .Y(n29) );
  NAND2X1 U31 ( .A(Cin), .B(n2), .Y(n33) );
  NAND2X1 U32 ( .A(n14), .B(n6), .Y(n66) );
  AND2X2 U33 ( .A(n55), .B(n52), .Y(n15) );
  OR2X2 U34 ( .A(B[2]), .B(A[2]), .Y(n53) );
  XOR2X1 U35 ( .A(n52), .B(n17), .Y(n63) );
  XNOR2X1 U36 ( .A(A[3]), .B(B[3]), .Y(n17) );
  XNOR2X1 U37 ( .A(Cin), .B(n18), .Y(S[0]) );
  XNOR2X1 U38 ( .A(B[0]), .B(n12), .Y(n18) );
  NAND2X1 U39 ( .A(n26), .B(n19), .Y(n54) );
  NAND2X1 U40 ( .A(n48), .B(n25), .Y(n21) );
  INVX2 U41 ( .A(B[0]), .Y(n28) );
  NOR2X1 U42 ( .A(n29), .B(n28), .Y(n23) );
  NAND2X1 U43 ( .A(A[1]), .B(B[1]), .Y(n36) );
  NAND2X1 U44 ( .A(A[2]), .B(B[2]), .Y(n52) );
  OAI21X1 U45 ( .A(n20), .B(n36), .C(n52), .Y(n22) );
  AOI22X1 U46 ( .A(PG), .B(n23), .C(n22), .D(n21), .Y(n24) );
  OAI21X1 U47 ( .A(n48), .B(n25), .C(n24), .Y(GG) );
  XOR2X1 U48 ( .A(n26), .B(A[1]), .Y(n32) );
  INVX2 U49 ( .A(n32), .Y(n27) );
  NAND2X1 U50 ( .A(B[0]), .B(A[0]), .Y(n37) );
  NAND2X1 U51 ( .A(n49), .B(n5), .Y(n35) );
  NAND2X1 U52 ( .A(n29), .B(n28), .Y(n56) );
  AOI22X1 U53 ( .A(n31), .B(n32), .C(n5), .D(n30), .Y(n34) );
  NAND3X1 U54 ( .A(n34), .B(n33), .C(n35), .Y(S[1]) );
  NAND2X1 U55 ( .A(n37), .B(n36), .Y(n38) );
  NAND2X1 U56 ( .A(n52), .B(n53), .Y(n43) );
  INVX2 U57 ( .A(n43), .Y(n44) );
  OAI21X1 U58 ( .A(n13), .B(n56), .C(n9), .Y(n39) );
  INVX2 U59 ( .A(n39), .Y(n42) );
  OAI21X1 U60 ( .A(n60), .B(n44), .C(n42), .Y(n41) );
  NAND2X1 U61 ( .A(n39), .B(n43), .Y(n40) );
  NAND2X1 U62 ( .A(n41), .B(n40), .Y(n47) );
  NAND3X1 U63 ( .A(n43), .B(Cin), .C(n42), .Y(n46) );
  NAND3X1 U64 ( .A(n47), .B(n46), .C(n45), .Y(S[2]) );
  XOR2X1 U65 ( .A(n48), .B(A[3]), .Y(n50) );
  INVX2 U66 ( .A(n50), .Y(n55) );
  NAND2X1 U67 ( .A(n16), .B(n50), .Y(n59) );
  NAND3X1 U68 ( .A(n55), .B(n9), .C(n53), .Y(n62) );
  NAND3X1 U69 ( .A(n57), .B(n60), .C(n15), .Y(n58) );
  OAI21X1 U70 ( .A(n60), .B(n59), .C(n58), .Y(n61) );
  NAND3X1 U71 ( .A(n64), .B(n65), .C(n66), .Y(S[3]) );
endmodule


module scalable_cla_block_CLA_BLK_SIZE_BITS4_1 ( A, B, Cin, S, PG, GG );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  INVX1 U1 ( .A(A[1]), .Y(n1) );
  INVX2 U2 ( .A(A[1]), .Y(n43) );
  INVX2 U3 ( .A(n50), .Y(n2) );
  INVX1 U4 ( .A(A[2]), .Y(n26) );
  INVX2 U5 ( .A(B[2]), .Y(n25) );
  BUFX2 U6 ( .A(n43), .Y(n3) );
  BUFX2 U7 ( .A(B[0]), .Y(n4) );
  AND2X2 U8 ( .A(n12), .B(n54), .Y(n5) );
  AND2X1 U9 ( .A(n51), .B(n52), .Y(n6) );
  INVX2 U10 ( .A(n57), .Y(n16) );
  XNOR2X1 U11 ( .A(n18), .B(n4), .Y(n7) );
  XNOR2X1 U12 ( .A(n22), .B(n7), .Y(S[0]) );
  BUFX2 U13 ( .A(n41), .Y(n8) );
  NAND2X1 U14 ( .A(n12), .B(n54), .Y(n9) );
  INVX1 U15 ( .A(n36), .Y(n37) );
  INVX2 U16 ( .A(n54), .Y(n20) );
  OR2X1 U17 ( .A(B[3]), .B(A[3]), .Y(n33) );
  BUFX2 U18 ( .A(B[3]), .Y(n17) );
  XNOR2X1 U19 ( .A(n17), .B(n50), .Y(n10) );
  INVX1 U20 ( .A(n10), .Y(n53) );
  INVX1 U21 ( .A(n16), .Y(n11) );
  INVX2 U22 ( .A(n14), .Y(n12) );
  INVX2 U23 ( .A(n59), .Y(n14) );
  INVX1 U24 ( .A(n42), .Y(n13) );
  NAND2X1 U25 ( .A(n22), .B(n6), .Y(n70) );
  INVX1 U26 ( .A(n64), .Y(n51) );
  INVX1 U27 ( .A(n14), .Y(n15) );
  INVX4 U28 ( .A(A[3]), .Y(n50) );
  BUFX2 U29 ( .A(A[0]), .Y(n18) );
  AND2X2 U30 ( .A(A[2]), .B(B[2]), .Y(n19) );
  INVX2 U31 ( .A(n19), .Y(n54) );
  INVX1 U32 ( .A(Cin), .Y(n66) );
  AND2X2 U33 ( .A(B[1]), .B(A[1]), .Y(n27) );
  OR2X2 U34 ( .A(n24), .B(B[3]), .Y(n21) );
  INVX2 U35 ( .A(n44), .Y(n46) );
  OR2X2 U36 ( .A(A[0]), .B(n4), .Y(n52) );
  BUFX4 U37 ( .A(Cin), .Y(n22) );
  INVX4 U38 ( .A(B[1]), .Y(n42) );
  INVX2 U39 ( .A(n50), .Y(n24) );
  OR2X1 U40 ( .A(n16), .B(n5), .Y(n23) );
  NAND2X1 U41 ( .A(n23), .B(n46), .Y(n45) );
  AOI22X1 U42 ( .A(n21), .B(n19), .C(n17), .D(n24), .Y(n32) );
  NAND2X1 U43 ( .A(n26), .B(n25), .Y(n59) );
  NAND3X1 U44 ( .A(n59), .B(n27), .C(n21), .Y(n31) );
  OAI21X1 U45 ( .A(B[3]), .B(n2), .C(B[0]), .Y(n28) );
  AOI21X1 U46 ( .A(n43), .B(n42), .C(n28), .Y(n29) );
  NAND3X1 U47 ( .A(A[0]), .B(n59), .C(n29), .Y(n30) );
  NAND3X1 U48 ( .A(n31), .B(n30), .C(n32), .Y(GG) );
  OAI21X1 U49 ( .A(A[2]), .B(B[2]), .C(n33), .Y(n34) );
  AOI21X1 U50 ( .A(n43), .B(n42), .C(n34), .Y(PG) );
  XOR2X1 U51 ( .A(n3), .B(n13), .Y(n36) );
  NAND3X1 U52 ( .A(n36), .B(n52), .C(n22), .Y(n40) );
  NAND2X1 U53 ( .A(B[0]), .B(A[0]), .Y(n41) );
  OAI21X1 U54 ( .A(n36), .B(n52), .C(n8), .Y(n35) );
  OAI21X1 U55 ( .A(n36), .B(n8), .C(n35), .Y(n39) );
  NAND3X1 U56 ( .A(n8), .B(n66), .C(n37), .Y(n38) );
  NAND3X1 U57 ( .A(n38), .B(n39), .C(n40), .Y(S[1]) );
  OAI21X1 U58 ( .A(n1), .B(n42), .C(n41), .Y(n57) );
  NAND3X1 U59 ( .A(n5), .B(n16), .C(n66), .Y(n49) );
  NAND2X1 U60 ( .A(n1), .B(n42), .Y(n60) );
  OAI21X1 U61 ( .A(n57), .B(n52), .C(n60), .Y(n44) );
  NAND3X1 U62 ( .A(n46), .B(n9), .C(n22), .Y(n48) );
  OAI21X1 U63 ( .A(n5), .B(n46), .C(n45), .Y(n47) );
  NAND3X1 U64 ( .A(n49), .B(n48), .C(n47), .Y(S[2]) );
  NAND3X1 U65 ( .A(n60), .B(n15), .C(n53), .Y(n64) );
  INVX2 U66 ( .A(n52), .Y(n56) );
  NAND2X1 U67 ( .A(n10), .B(n54), .Y(n58) );
  INVX2 U68 ( .A(n58), .Y(n55) );
  NAND3X1 U69 ( .A(n56), .B(n16), .C(n55), .Y(n69) );
  NOR2X1 U70 ( .A(n58), .B(n11), .Y(n67) );
  NAND2X1 U71 ( .A(n60), .B(n10), .Y(n62) );
  XOR2X1 U72 ( .A(n10), .B(n20), .Y(n61) );
  OAI21X1 U73 ( .A(n14), .B(n62), .C(n61), .Y(n63) );
  OAI21X1 U74 ( .A(n16), .B(n64), .C(n63), .Y(n65) );
  AOI21X1 U75 ( .A(n67), .B(n66), .C(n65), .Y(n68) );
  NAND3X1 U76 ( .A(n69), .B(n70), .C(n68), .Y(S[3]) );
endmodule


module scalable_cla_block_CLA_BLK_SIZE_BITS4_2 ( A, B, Cin, S, PG, GG );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  output PG, GG;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;

  INVX1 U1 ( .A(n41), .Y(n1) );
  OR2X2 U2 ( .A(n7), .B(n2), .Y(n35) );
  INVX2 U3 ( .A(B[3]), .Y(n39) );
  BUFX2 U4 ( .A(A[0]), .Y(n2) );
  INVX2 U5 ( .A(B[2]), .Y(n12) );
  INVX2 U6 ( .A(A[3]), .Y(n22) );
  XOR2X1 U7 ( .A(n3), .B(n19), .Y(S[0]) );
  INVX1 U8 ( .A(n1), .Y(n3) );
  XOR2X1 U9 ( .A(n4), .B(n2), .Y(n19) );
  INVX1 U10 ( .A(n7), .Y(n4) );
  XNOR2X1 U11 ( .A(n38), .B(n5), .Y(S[2]) );
  OR2X2 U12 ( .A(n49), .B(n43), .Y(n5) );
  BUFX2 U13 ( .A(n39), .Y(n6) );
  BUFX2 U14 ( .A(B[0]), .Y(n7) );
  BUFX2 U15 ( .A(n46), .Y(n8) );
  INVX1 U16 ( .A(n34), .Y(n9) );
  INVX1 U17 ( .A(n23), .Y(n43) );
  INVX2 U18 ( .A(n15), .Y(n10) );
  INVX1 U19 ( .A(n39), .Y(n11) );
  NAND2X1 U20 ( .A(n12), .B(n13), .Y(n14) );
  NAND2X1 U21 ( .A(n14), .B(B[1]), .Y(n21) );
  INVX1 U22 ( .A(A[2]), .Y(n13) );
  BUFX2 U23 ( .A(n33), .Y(n15) );
  OR2X2 U24 ( .A(B[1]), .B(A[1]), .Y(n46) );
  INVX1 U25 ( .A(n22), .Y(n16) );
  INVX2 U26 ( .A(B[3]), .Y(n17) );
  NAND2X1 U27 ( .A(n33), .B(n34), .Y(n18) );
  OR2X2 U28 ( .A(A[2]), .B(B[2]), .Y(n44) );
  XNOR2X1 U29 ( .A(n31), .B(n20), .Y(S[1]) );
  XNOR2X1 U30 ( .A(n10), .B(n9), .Y(n20) );
  NAND2X1 U31 ( .A(n39), .B(n22), .Y(n29) );
  INVX2 U32 ( .A(B[1]), .Y(n34) );
  INVX2 U33 ( .A(A[1]), .Y(n33) );
  NAND2X1 U34 ( .A(n18), .B(n29), .Y(n28) );
  NAND3X1 U35 ( .A(n44), .B(A[0]), .C(B[0]), .Y(n27) );
  NAND2X1 U36 ( .A(B[2]), .B(A[2]), .Y(n23) );
  AOI22X1 U37 ( .A(n22), .B(n17), .C(n23), .D(n21), .Y(n25) );
  NAND2X1 U38 ( .A(n23), .B(n33), .Y(n24) );
  AOI22X1 U39 ( .A(n24), .B(n25), .C(A[3]), .D(n11), .Y(n26) );
  OAI21X1 U40 ( .A(n28), .B(n27), .C(n26), .Y(GG) );
  NAND3X1 U41 ( .A(n44), .B(n46), .C(n29), .Y(n30) );
  INVX2 U42 ( .A(n30), .Y(PG) );
  INVX2 U43 ( .A(n35), .Y(n42) );
  INVX2 U44 ( .A(Cin), .Y(n41) );
  NAND2X1 U45 ( .A(A[0]), .B(B[0]), .Y(n32) );
  OAI21X1 U46 ( .A(n41), .B(n42), .C(n32), .Y(n31) );
  OAI21X1 U47 ( .A(n34), .B(n15), .C(n32), .Y(n36) );
  INVX2 U48 ( .A(n36), .Y(n40) );
  OAI21X1 U49 ( .A(n36), .B(n35), .C(n8), .Y(n37) );
  AOI21X1 U50 ( .A(n41), .B(n40), .C(n37), .Y(n38) );
  INVX2 U51 ( .A(n44), .Y(n49) );
  XOR2X1 U52 ( .A(n6), .B(n16), .Y(n47) );
  INVX2 U53 ( .A(n47), .Y(n45) );
  NAND2X1 U54 ( .A(n23), .B(n45), .Y(n55) );
  OAI21X1 U55 ( .A(n41), .B(n42), .C(n40), .Y(n54) );
  XOR2X1 U56 ( .A(n45), .B(n43), .Y(n52) );
  NAND3X1 U57 ( .A(n45), .B(n18), .C(n44), .Y(n51) );
  NAND2X1 U58 ( .A(n47), .B(n8), .Y(n48) );
  NOR2X1 U59 ( .A(n49), .B(n48), .Y(n50) );
  AOI22X1 U60 ( .A(n52), .B(n51), .C(n54), .D(n50), .Y(n53) );
  OAI21X1 U61 ( .A(n54), .B(n55), .C(n53), .Y(S[3]) );
endmodule


module scalable_cla_addr_NUM_CLA_BLKS4_CLA_BLK_SIZE_BITS4 ( A, B, Cin, S, V );
  input [15:0] A;
  input [15:0] B;
  output [15:0] S;
  input Cin;
  output V;
  wire   n2, n3, n4, n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [3:0] gg_vector;
  wire   [3:0] pg_vector;

  scalable_cla_block_CLA_BLK_SIZE_BITS4_3 CLA_BLK_0 ( .A(A[3:0]), .B(B[3:0]), 
        .Cin(Cin), .S(S[3:0]), .PG(pg_vector[0]), .GG(gg_vector[0]) );
  scalable_cla_block_CLA_BLK_SIZE_BITS4_2 CLA_BLK_1 ( .A(A[7:4]), .B(B[7:4]), 
        .Cin(n4), .S(S[7:4]), .PG(pg_vector[1]), .GG(gg_vector[1]) );
  scalable_cla_block_CLA_BLK_SIZE_BITS4_1 CLA_BLK_2 ( .A(A[11:8]), .B(B[11:8]), 
        .Cin(n3), .S(S[11:8]), .PG(pg_vector[2]), .GG(gg_vector[2]) );
  scalable_cla_block_CLA_BLK_SIZE_BITS4_0 CLA_BLK_3 ( .A(A[15:12]), .B(
        B[15:12]), .Cin(n1), .S(S[15:12]), .PG(pg_vector[3]), .GG(gg_vector[3]) );
  INVX1 U1 ( .A(n14), .Y(V) );
  BUFX4 U2 ( .A(n2), .Y(n1) );
  BUFX2 U3 ( .A(n1), .Y(n5) );
  INVX1 U4 ( .A(gg_vector[0]), .Y(n13) );
  INVX1 U5 ( .A(gg_vector[1]), .Y(n11) );
  NAND2X1 U6 ( .A(pg_vector[0]), .B(Cin), .Y(n12) );
  INVX2 U7 ( .A(n12), .Y(n9) );
  NOR2X1 U8 ( .A(n9), .B(gg_vector[0]), .Y(n8) );
  NAND2X1 U9 ( .A(pg_vector[1]), .B(pg_vector[2]), .Y(n7) );
  AOI21X1 U10 ( .A(pg_vector[2]), .B(gg_vector[1]), .C(gg_vector[2]), .Y(n6)
         );
  OAI21X1 U11 ( .A(n7), .B(n8), .C(n6), .Y(n2) );
  OAI21X1 U12 ( .A(gg_vector[0]), .B(n9), .C(pg_vector[1]), .Y(n10) );
  NAND2X1 U13 ( .A(n10), .B(n11), .Y(n3) );
  NAND2X1 U14 ( .A(n12), .B(n13), .Y(n4) );
  AOI21X1 U15 ( .A(pg_vector[3]), .B(n5), .C(gg_vector[3]), .Y(n14) );
endmodule


module alu_DATA_SIZE_BITS16 ( A, B, alu_op, result, overflow );
  input [15:0] A;
  input [15:0] B;
  output [15:0] result;
  input alu_op;
  output overflow;
  wire   int_V, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50;
  wire   [15:0] int_A;
  wire   [15:0] int_B;
  wire   [15:0] int_S;

  scalable_cla_addr_NUM_CLA_BLKS4_CLA_BLK_SIZE_BITS4 CLA_ADDR ( .A(int_A), .B(
        int_B), .Cin(1'b0), .S(int_S), .V(int_V) );
  AND2X2 U2 ( .A(alu_op), .B(A[14]), .Y(int_A[14]) );
  INVX1 U3 ( .A(A[14]), .Y(n34) );
  INVX1 U4 ( .A(n26), .Y(n22) );
  INVX2 U5 ( .A(n26), .Y(n3) );
  MUX2X1 U6 ( .B(n4), .A(int_S[14]), .S(n8), .Y(n49) );
  BUFX2 U7 ( .A(A[3]), .Y(n1) );
  INVX1 U8 ( .A(n33), .Y(n2) );
  AND2X2 U9 ( .A(n3), .B(A[6]), .Y(int_A[6]) );
  INVX1 U10 ( .A(A[6]), .Y(n31) );
  INVX1 U11 ( .A(n39), .Y(result[4]) );
  INVX1 U12 ( .A(n34), .Y(n4) );
  INVX1 U13 ( .A(n43), .Y(result[8]) );
  INVX1 U14 ( .A(n47), .Y(result[12]) );
  INVX1 U15 ( .A(n31), .Y(n5) );
  INVX1 U16 ( .A(n49), .Y(result[14]) );
  INVX1 U17 ( .A(n50), .Y(result[15]) );
  AND2X2 U18 ( .A(A[10]), .B(alu_op), .Y(int_A[10]) );
  INVX1 U19 ( .A(A[10]), .Y(n32) );
  BUFX2 U20 ( .A(A[7]), .Y(n6) );
  AND2X2 U21 ( .A(n25), .B(A[1]), .Y(int_A[1]) );
  INVX1 U22 ( .A(A[1]), .Y(n27) );
  INVX1 U23 ( .A(n30), .Y(n7) );
  AND2X2 U24 ( .A(n25), .B(A[2]), .Y(int_A[2]) );
  INVX4 U25 ( .A(n26), .Y(n8) );
  BUFX2 U26 ( .A(A[0]), .Y(n9) );
  INVX1 U27 ( .A(n29), .Y(n10) );
  BUFX2 U28 ( .A(A[9]), .Y(n11) );
  INVX1 U29 ( .A(n27), .Y(n12) );
  INVX2 U30 ( .A(n26), .Y(n13) );
  NAND2X1 U31 ( .A(n13), .B(A[7]), .Y(n14) );
  INVX2 U32 ( .A(n14), .Y(int_A[7]) );
  INVX2 U33 ( .A(n26), .Y(n25) );
  AND2X2 U34 ( .A(A[15]), .B(n13), .Y(int_A[15]) );
  BUFX2 U35 ( .A(A[11]), .Y(n15) );
  INVX8 U36 ( .A(alu_op), .Y(n26) );
  INVX1 U37 ( .A(n44), .Y(result[9]) );
  INVX2 U38 ( .A(n26), .Y(n24) );
  INVX2 U39 ( .A(A[5]), .Y(n30) );
  INVX2 U40 ( .A(n26), .Y(n21) );
  INVX2 U41 ( .A(n13), .Y(n16) );
  INVX4 U42 ( .A(n16), .Y(n17) );
  INVX1 U43 ( .A(A[2]), .Y(n28) );
  INVX1 U44 ( .A(n41), .Y(result[6]) );
  INVX1 U45 ( .A(n32), .Y(n18) );
  INVX1 U46 ( .A(n28), .Y(n19) );
  INVX1 U47 ( .A(n40), .Y(result[5]) );
  INVX1 U48 ( .A(n26), .Y(n20) );
  AND2X1 U49 ( .A(A[15]), .B(n26), .Y(n23) );
  AND2X2 U50 ( .A(n20), .B(A[3]), .Y(int_A[3]) );
  AND2X2 U51 ( .A(n21), .B(A[13]), .Y(int_A[13]) );
  AND2X2 U52 ( .A(n22), .B(A[11]), .Y(int_A[11]) );
  AND2X2 U53 ( .A(A[9]), .B(n17), .Y(int_A[9]) );
  INVX1 U54 ( .A(n48), .Y(result[13]) );
  AND2X2 U55 ( .A(n8), .B(A[8]), .Y(int_A[8]) );
  INVX1 U56 ( .A(n42), .Y(result[7]) );
  INVX1 U57 ( .A(n46), .Y(result[11]) );
  INVX1 U58 ( .A(n45), .Y(result[10]) );
  AND2X2 U59 ( .A(n24), .B(A[0]), .Y(int_A[0]) );
  AND2X2 U60 ( .A(B[0]), .B(n13), .Y(int_B[0]) );
  AND2X2 U61 ( .A(B[1]), .B(n3), .Y(int_B[1]) );
  AND2X2 U62 ( .A(n25), .B(B[2]), .Y(int_B[2]) );
  AND2X2 U63 ( .A(n25), .B(B[3]), .Y(int_B[3]) );
  AND2X2 U64 ( .A(B[4]), .B(n24), .Y(int_B[4]) );
  AND2X2 U65 ( .A(B[5]), .B(n20), .Y(int_B[5]) );
  AND2X2 U66 ( .A(B[6]), .B(n22), .Y(int_B[6]) );
  AND2X2 U67 ( .A(n21), .B(B[7]), .Y(int_B[7]) );
  AND2X2 U68 ( .A(B[8]), .B(n21), .Y(int_B[8]) );
  AND2X2 U69 ( .A(B[9]), .B(n17), .Y(int_B[9]) );
  AND2X2 U70 ( .A(B[10]), .B(n24), .Y(int_B[10]) );
  AND2X2 U71 ( .A(B[11]), .B(n3), .Y(int_B[11]) );
  AND2X2 U72 ( .A(B[12]), .B(n8), .Y(int_B[12]) );
  AND2X2 U73 ( .A(B[13]), .B(n24), .Y(int_B[13]) );
  AND2X2 U74 ( .A(B[14]), .B(n17), .Y(int_B[14]) );
  AND2X2 U75 ( .A(B[15]), .B(n21), .Y(int_B[15]) );
  INVX2 U76 ( .A(A[4]), .Y(n29) );
  NOR2X1 U77 ( .A(n26), .B(n29), .Y(int_A[4]) );
  NOR2X1 U78 ( .A(n26), .B(n30), .Y(int_A[5]) );
  INVX2 U79 ( .A(A[12]), .Y(n33) );
  NOR2X1 U80 ( .A(n26), .B(n33), .Y(int_A[12]) );
  AND2X2 U81 ( .A(int_V), .B(n8), .Y(overflow) );
  MUX2X1 U82 ( .B(n9), .A(int_S[0]), .S(n8), .Y(n35) );
  INVX2 U83 ( .A(n35), .Y(result[0]) );
  MUX2X1 U84 ( .B(n12), .A(int_S[1]), .S(n8), .Y(n36) );
  INVX2 U85 ( .A(n36), .Y(result[1]) );
  MUX2X1 U86 ( .B(n19), .A(int_S[2]), .S(n8), .Y(n37) );
  INVX2 U87 ( .A(n37), .Y(result[2]) );
  MUX2X1 U88 ( .B(n1), .A(int_S[3]), .S(n8), .Y(n38) );
  INVX2 U89 ( .A(n38), .Y(result[3]) );
  MUX2X1 U90 ( .B(n10), .A(int_S[4]), .S(n8), .Y(n39) );
  MUX2X1 U91 ( .B(n7), .A(int_S[5]), .S(n8), .Y(n40) );
  MUX2X1 U92 ( .B(n5), .A(int_S[6]), .S(n8), .Y(n41) );
  MUX2X1 U93 ( .B(n6), .A(int_S[7]), .S(n8), .Y(n42) );
  MUX2X1 U94 ( .B(A[8]), .A(int_S[8]), .S(n8), .Y(n43) );
  MUX2X1 U95 ( .B(n11), .A(int_S[9]), .S(n8), .Y(n44) );
  MUX2X1 U96 ( .B(n18), .A(int_S[10]), .S(n8), .Y(n45) );
  MUX2X1 U97 ( .B(n15), .A(int_S[11]), .S(n8), .Y(n46) );
  MUX2X1 U98 ( .B(n2), .A(int_S[12]), .S(n8), .Y(n47) );
  MUX2X1 U99 ( .B(A[13]), .A(int_S[13]), .S(n8), .Y(n48) );
  OAI22X1 U100 ( .A(n17), .B(n23), .C(n23), .D(int_S[15]), .Y(n50) );
endmodule


module datapath ( clk, n_reset, op, src1, src2, dest, ext_data, outreg_data, 
        overflow );
  input [1:0] op;
  input [3:0] src1;
  input [3:0] src2;
  input [3:0] dest;
  input [15:0] ext_data;
  output [15:0] outreg_data;
  input clk, n_reset;
  output overflow;
  wire   int_w_data_sel, int_w_en, int_alu_op, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  wire   [15:0] int_src1_data;
  wire   [15:0] int_src2_data;
  wire   [15:0] int_result;

  datapath_ctrl DP_CTRL ( .op(op), .w_data_sel(int_w_data_sel), .w_en(int_w_en), .alu_op(int_alu_op) );
  regfile_NUM_REG_ADDR_BITS4_REG_SIZE_BITS16 REG_FILE ( .clk(clk), .n_reset(
        n_reset), .w_sel(dest), .r1_sel(src1), .r2_sel(src2), .w_data({n10, 
        n11, n12, n13, n14, n15, n1, n2, n3, n4, n5, n6, n7, n8, n9, n16}), 
        .w_en(int_w_en), .r1_data(int_src1_data), .r2_data(int_src2_data), 
        .outreg_data(outreg_data) );
  alu_DATA_SIZE_BITS16 ALU_MAP ( .A(int_src1_data), .B(int_src2_data), 
        .alu_op(int_alu_op), .result(int_result), .overflow(overflow) );
  INVX4 U1 ( .A(n21), .Y(n9) );
  INVX4 U2 ( .A(n24), .Y(n6) );
  INVX4 U3 ( .A(n23), .Y(n7) );
  INVX4 U4 ( .A(n22), .Y(n8) );
  INVX4 U5 ( .A(n28), .Y(n2) );
  INVX4 U6 ( .A(n25), .Y(n5) );
  INVX2 U7 ( .A(n18), .Y(n35) );
  INVX2 U8 ( .A(n17), .Y(n18) );
  INVX2 U9 ( .A(n17), .Y(n19) );
  INVX1 U10 ( .A(int_w_data_sel), .Y(n17) );
  INVX4 U11 ( .A(n26), .Y(n4) );
  INVX4 U12 ( .A(n32), .Y(n13) );
  INVX4 U13 ( .A(n27), .Y(n3) );
  INVX4 U14 ( .A(n29), .Y(n1) );
  INVX4 U15 ( .A(n34), .Y(n11) );
  INVX4 U16 ( .A(n36), .Y(n10) );
  INVX4 U17 ( .A(n31), .Y(n14) );
  INVX4 U18 ( .A(n33), .Y(n12) );
  INVX4 U19 ( .A(n30), .Y(n15) );
  MUX2X1 U20 ( .B(ext_data[0]), .A(int_result[0]), .S(n18), .Y(n20) );
  INVX2 U21 ( .A(n20), .Y(n16) );
  MUX2X1 U22 ( .B(ext_data[1]), .A(int_result[1]), .S(n18), .Y(n21) );
  MUX2X1 U23 ( .B(ext_data[2]), .A(int_result[2]), .S(n18), .Y(n22) );
  MUX2X1 U24 ( .B(ext_data[3]), .A(int_result[3]), .S(n18), .Y(n23) );
  MUX2X1 U25 ( .B(ext_data[4]), .A(int_result[4]), .S(n18), .Y(n24) );
  AOI22X1 U26 ( .A(int_result[5]), .B(n19), .C(ext_data[5]), .D(n35), .Y(n25)
         );
  AOI22X1 U27 ( .A(int_result[6]), .B(n19), .C(ext_data[6]), .D(n35), .Y(n26)
         );
  AOI22X1 U28 ( .A(int_result[7]), .B(n19), .C(ext_data[7]), .D(n35), .Y(n27)
         );
  AOI22X1 U29 ( .A(int_result[8]), .B(n19), .C(ext_data[8]), .D(n35), .Y(n28)
         );
  AOI22X1 U30 ( .A(int_result[9]), .B(n19), .C(ext_data[9]), .D(n35), .Y(n29)
         );
  AOI22X1 U31 ( .A(int_result[10]), .B(n19), .C(ext_data[10]), .D(n35), .Y(n30) );
  AOI22X1 U32 ( .A(int_result[11]), .B(n19), .C(ext_data[11]), .D(n35), .Y(n31) );
  AOI22X1 U33 ( .A(int_result[12]), .B(n19), .C(ext_data[12]), .D(n35), .Y(n32) );
  AOI22X1 U34 ( .A(int_result[13]), .B(n19), .C(ext_data[13]), .D(n35), .Y(n33) );
  AOI22X1 U35 ( .A(ext_data[14]), .B(n35), .C(int_result[14]), .D(n18), .Y(n34) );
  AOI22X1 U36 ( .A(ext_data[15]), .B(n35), .C(int_result[15]), .D(n19), .Y(n36) );
endmodule


module counter ( clk, n_reset, cnt_up, one_k_samples );
  input clk, n_reset, cnt_up;
  output one_k_samples;
  wire   nextflag, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n18, n20, n22;
  wire   [3:0] counter;

  DFFSR \counter_reg[0]  ( .D(n22), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        counter[0]) );
  DFFSR \counter_reg[1]  ( .D(n20), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        counter[1]) );
  DFFSR \counter_reg[2]  ( .D(n18), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        counter[2]) );
  DFFSR \counter_reg[3]  ( .D(n16), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        counter[3]) );
  DFFSR flagger_reg ( .D(nextflag), .CLK(clk), .R(n_reset), .S(1'b1), .Q(
        one_k_samples) );
  NOR2X1 U3 ( .A(n5), .B(n6), .Y(nextflag) );
  XNOR2X1 U4 ( .A(counter[3]), .B(n6), .Y(n16) );
  NAND2X1 U5 ( .A(counter[2]), .B(n7), .Y(n6) );
  XOR2X1 U6 ( .A(counter[2]), .B(n7), .Y(n18) );
  NOR2X1 U7 ( .A(n8), .B(n9), .Y(n7) );
  INVX1 U8 ( .A(counter[1]), .Y(n8) );
  XNOR2X1 U9 ( .A(counter[1]), .B(n9), .Y(n20) );
  NAND2X1 U10 ( .A(counter[0]), .B(cnt_up), .Y(n9) );
  OAI21X1 U11 ( .A(counter[0]), .B(n10), .C(n11), .Y(n22) );
  NAND2X1 U12 ( .A(counter[0]), .B(n12), .Y(n11) );
  OAI21X1 U13 ( .A(n5), .B(n13), .C(cnt_up), .Y(n12) );
  NAND2X1 U14 ( .A(counter[2]), .B(counter[1]), .Y(n13) );
  INVX1 U15 ( .A(counter[3]), .Y(n5) );
  INVX1 U16 ( .A(cnt_up), .Y(n10) );
endmodule


module avg_four ( clk, n_reset, sample_data, data_ready, one_k_samples, 
        modwait, avg_out, err );
  input [15:0] sample_data;
  output [15:0] avg_out;
  input clk, n_reset, data_ready;
  output one_k_samples, modwait, err;
  wire   dr, test_overflow, count_en;
  wire   [1:0] op;
  wire   [3:0] src1;
  wire   [3:0] src2;
  wire   [3:0] dest;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign avg_out[14] = 1'b0;
  assign avg_out[15] = 1'b0;

  sync U2 ( .clk(clk), .n_reset(n_reset), .async_in(data_ready), .sync_out(dr)
         );
  controller U1 ( .clk(clk), .n_reset(n_reset), .dr(dr), .overflow(
        test_overflow), .cnt_up(count_en), .modwait(modwait), .op(op), .src1(
        src1), .src2(src2), .dest(dest), .err(err) );
  datapath U3 ( .clk(clk), .n_reset(n_reset), .op(op), .src1({1'b0, src1[2:0]}), .src2({1'b0, src2[2:0]}), .dest({1'b0, dest[2:0]}), .ext_data(sample_data), 
        .outreg_data({avg_out[13:0], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}), .overflow(test_overflow) );
  counter U4 ( .clk(clk), .n_reset(n_reset), .cnt_up(count_en), 
        .one_k_samples(one_k_samples) );
endmodule

